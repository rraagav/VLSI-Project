magic
tech scmos
timestamp 1700503255
<< nwell >>
rect 71 48 131 72
rect 669 48 729 72
rect 1548 48 1608 72
rect 2316 48 2376 72
rect -2 0 58 24
rect 172 -20 232 4
rect 596 0 656 24
rect 770 -20 830 4
rect 1475 0 1535 24
rect 1649 -20 1709 4
rect 2243 0 2303 24
rect 2417 -20 2477 4
rect 86 -61 146 -37
rect 684 -61 744 -37
rect 1563 -61 1623 -37
rect 2331 -61 2391 -37
rect 352 -255 412 -231
rect 1095 -258 1155 -234
rect 1854 -258 1914 -234
rect 2590 -258 2650 -234
rect 42 -303 102 -279
rect 279 -303 339 -279
rect 453 -323 513 -299
rect 785 -306 845 -282
rect 1022 -306 1082 -282
rect 1196 -326 1256 -302
rect 1544 -306 1604 -282
rect 1781 -306 1841 -282
rect 1955 -326 2015 -302
rect 2280 -306 2340 -282
rect 2517 -306 2577 -282
rect 2691 -326 2751 -302
rect -31 -351 29 -327
rect 143 -371 203 -347
rect 367 -364 427 -340
rect 712 -354 772 -330
rect 886 -374 946 -350
rect 1110 -367 1170 -343
rect 1471 -354 1531 -330
rect 1645 -374 1705 -350
rect 1869 -367 1929 -343
rect 2207 -354 2267 -330
rect 2381 -374 2441 -350
rect 2605 -367 2665 -343
rect 57 -412 117 -388
rect 800 -415 860 -391
rect 1559 -415 1619 -391
rect 2295 -415 2355 -391
rect 339 -470 399 -446
rect 405 -470 433 -446
rect 498 -470 558 -446
rect 566 -470 594 -446
rect 1082 -473 1142 -449
rect 1148 -473 1176 -449
rect 1241 -473 1301 -449
rect 1309 -473 1337 -449
rect 1841 -473 1901 -449
rect 1907 -473 1935 -449
rect 2000 -473 2060 -449
rect 2068 -473 2096 -449
rect 2577 -473 2637 -449
rect 2643 -473 2671 -449
rect 2736 -473 2796 -449
rect 2804 -473 2832 -449
rect 28 -521 88 -497
rect 94 -521 122 -497
rect 771 -524 831 -500
rect 837 -524 865 -500
rect 1530 -524 1590 -500
rect 1596 -524 1624 -500
rect 2266 -524 2326 -500
rect 2332 -524 2360 -500
<< ntransistor >>
rect 83 11 87 19
rect 104 11 108 19
rect 681 11 685 19
rect 702 11 706 19
rect 10 -37 14 -29
rect 31 -37 35 -29
rect 1560 11 1564 19
rect 1581 11 1585 19
rect 608 -37 612 -29
rect 629 -37 633 -29
rect 184 -57 188 -49
rect 205 -57 209 -49
rect 2328 11 2332 19
rect 2349 11 2353 19
rect 1487 -37 1491 -29
rect 1508 -37 1512 -29
rect 782 -57 786 -49
rect 803 -57 807 -49
rect 2255 -37 2259 -29
rect 2276 -37 2280 -29
rect 1661 -57 1665 -49
rect 1682 -57 1686 -49
rect 2429 -57 2433 -49
rect 2450 -57 2454 -49
rect 98 -98 102 -90
rect 119 -98 123 -90
rect 696 -98 700 -90
rect 717 -98 721 -90
rect 1575 -98 1579 -90
rect 1596 -98 1600 -90
rect 2343 -98 2347 -90
rect 2364 -98 2368 -90
rect 364 -292 368 -284
rect 385 -292 389 -284
rect 1107 -295 1111 -287
rect 1128 -295 1132 -287
rect 54 -340 58 -332
rect 75 -340 79 -332
rect 291 -340 295 -332
rect 312 -340 316 -332
rect 1866 -295 1870 -287
rect 1887 -295 1891 -287
rect 797 -343 801 -335
rect 818 -343 822 -335
rect 1034 -343 1038 -335
rect 1055 -343 1059 -335
rect -19 -388 -15 -380
rect 2 -388 6 -380
rect 465 -360 469 -352
rect 486 -360 490 -352
rect 2602 -295 2606 -287
rect 2623 -295 2627 -287
rect 1556 -343 1560 -335
rect 1577 -343 1581 -335
rect 1793 -343 1797 -335
rect 1814 -343 1818 -335
rect 724 -391 728 -383
rect 745 -391 749 -383
rect 155 -408 159 -400
rect 176 -408 180 -400
rect 379 -401 383 -393
rect 400 -401 404 -393
rect 1208 -363 1212 -355
rect 1229 -363 1233 -355
rect 2292 -343 2296 -335
rect 2313 -343 2317 -335
rect 2529 -343 2533 -335
rect 2550 -343 2554 -335
rect 1483 -391 1487 -383
rect 1504 -391 1508 -383
rect 69 -449 73 -441
rect 90 -449 94 -441
rect 898 -411 902 -403
rect 919 -411 923 -403
rect 1122 -404 1126 -396
rect 1143 -404 1147 -396
rect 1967 -363 1971 -355
rect 1988 -363 1992 -355
rect 2219 -391 2223 -383
rect 2240 -391 2244 -383
rect 1657 -411 1661 -403
rect 1678 -411 1682 -403
rect 1881 -404 1885 -396
rect 1902 -404 1906 -396
rect 2703 -363 2707 -355
rect 2724 -363 2728 -355
rect 2393 -411 2397 -403
rect 2414 -411 2418 -403
rect 2617 -404 2621 -396
rect 2638 -404 2642 -396
rect 812 -452 816 -444
rect 833 -452 837 -444
rect 1571 -452 1575 -444
rect 1592 -452 1596 -444
rect 2307 -452 2311 -444
rect 2328 -452 2332 -444
rect 351 -507 355 -499
rect 372 -507 376 -499
rect 417 -507 421 -499
rect 510 -510 514 -502
rect 531 -510 535 -502
rect 578 -510 582 -502
rect 1094 -510 1098 -502
rect 1115 -510 1119 -502
rect 1160 -510 1164 -502
rect 1253 -513 1257 -505
rect 1274 -513 1278 -505
rect 1321 -513 1325 -505
rect 1853 -510 1857 -502
rect 1874 -510 1878 -502
rect 1919 -510 1923 -502
rect 2012 -513 2016 -505
rect 2033 -513 2037 -505
rect 2080 -513 2084 -505
rect 2589 -510 2593 -502
rect 2610 -510 2614 -502
rect 2655 -510 2659 -502
rect 2748 -513 2752 -505
rect 2769 -513 2773 -505
rect 2816 -513 2820 -505
rect 40 -558 44 -550
rect 61 -558 65 -550
rect 106 -558 110 -550
rect 783 -561 787 -553
rect 804 -561 808 -553
rect 849 -561 853 -553
rect 1542 -561 1546 -553
rect 1563 -561 1567 -553
rect 1608 -561 1612 -553
rect 2278 -561 2282 -553
rect 2299 -561 2303 -553
rect 2344 -561 2348 -553
<< ptransistor >>
rect 83 56 87 64
rect 104 56 108 64
rect 681 56 685 64
rect 702 56 706 64
rect 1560 56 1564 64
rect 1581 56 1585 64
rect 2328 56 2332 64
rect 2349 56 2353 64
rect 10 8 14 16
rect 31 8 35 16
rect 608 8 612 16
rect 629 8 633 16
rect 184 -12 188 -4
rect 205 -12 209 -4
rect 98 -53 102 -45
rect 119 -53 123 -45
rect 1487 8 1491 16
rect 1508 8 1512 16
rect 782 -12 786 -4
rect 803 -12 807 -4
rect 696 -53 700 -45
rect 717 -53 721 -45
rect 2255 8 2259 16
rect 2276 8 2280 16
rect 1661 -12 1665 -4
rect 1682 -12 1686 -4
rect 1575 -53 1579 -45
rect 1596 -53 1600 -45
rect 2429 -12 2433 -4
rect 2450 -12 2454 -4
rect 2343 -53 2347 -45
rect 2364 -53 2368 -45
rect 364 -247 368 -239
rect 385 -247 389 -239
rect 1107 -250 1111 -242
rect 1128 -250 1132 -242
rect 1866 -250 1870 -242
rect 1887 -250 1891 -242
rect 2602 -250 2606 -242
rect 2623 -250 2627 -242
rect 54 -295 58 -287
rect 75 -295 79 -287
rect 291 -295 295 -287
rect 312 -295 316 -287
rect 797 -298 801 -290
rect 818 -298 822 -290
rect 1034 -298 1038 -290
rect 1055 -298 1059 -290
rect 465 -315 469 -307
rect 486 -315 490 -307
rect -19 -343 -15 -335
rect 2 -343 6 -335
rect 155 -363 159 -355
rect 176 -363 180 -355
rect 379 -356 383 -348
rect 400 -356 404 -348
rect 1556 -298 1560 -290
rect 1577 -298 1581 -290
rect 1793 -298 1797 -290
rect 1814 -298 1818 -290
rect 1208 -318 1212 -310
rect 1229 -318 1233 -310
rect 724 -346 728 -338
rect 745 -346 749 -338
rect 69 -404 73 -396
rect 90 -404 94 -396
rect 898 -366 902 -358
rect 919 -366 923 -358
rect 1122 -359 1126 -351
rect 1143 -359 1147 -351
rect 2292 -298 2296 -290
rect 2313 -298 2317 -290
rect 2529 -298 2533 -290
rect 2550 -298 2554 -290
rect 1967 -318 1971 -310
rect 1988 -318 1992 -310
rect 1483 -346 1487 -338
rect 1504 -346 1508 -338
rect 812 -407 816 -399
rect 833 -407 837 -399
rect 1657 -366 1661 -358
rect 1678 -366 1682 -358
rect 1881 -359 1885 -351
rect 1902 -359 1906 -351
rect 2703 -318 2707 -310
rect 2724 -318 2728 -310
rect 2219 -346 2223 -338
rect 2240 -346 2244 -338
rect 1571 -407 1575 -399
rect 1592 -407 1596 -399
rect 2393 -366 2397 -358
rect 2414 -366 2418 -358
rect 2617 -359 2621 -351
rect 2638 -359 2642 -351
rect 2307 -407 2311 -399
rect 2328 -407 2332 -399
rect 351 -462 355 -454
rect 372 -462 376 -454
rect 417 -462 421 -454
rect 510 -462 514 -454
rect 531 -462 535 -454
rect 578 -462 582 -454
rect 40 -513 44 -505
rect 61 -513 65 -505
rect 106 -513 110 -505
rect 1094 -465 1098 -457
rect 1115 -465 1119 -457
rect 1160 -465 1164 -457
rect 1253 -465 1257 -457
rect 1274 -465 1278 -457
rect 1321 -465 1325 -457
rect 1853 -465 1857 -457
rect 1874 -465 1878 -457
rect 1919 -465 1923 -457
rect 2012 -465 2016 -457
rect 2033 -465 2037 -457
rect 2080 -465 2084 -457
rect 2589 -465 2593 -457
rect 2610 -465 2614 -457
rect 2655 -465 2659 -457
rect 2748 -465 2752 -457
rect 2769 -465 2773 -457
rect 2816 -465 2820 -457
rect 783 -516 787 -508
rect 804 -516 808 -508
rect 849 -516 853 -508
rect 1542 -516 1546 -508
rect 1563 -516 1567 -508
rect 1608 -516 1612 -508
rect 2278 -516 2282 -508
rect 2299 -516 2303 -508
rect 2344 -516 2348 -508
<< ndiffusion >>
rect 77 17 83 19
rect 77 13 78 17
rect 82 13 83 17
rect 77 11 83 13
rect 87 11 104 19
rect 108 17 125 19
rect 108 13 111 17
rect 115 13 125 17
rect 675 17 681 19
rect 108 11 125 13
rect 675 13 676 17
rect 680 13 681 17
rect 675 11 681 13
rect 685 11 702 19
rect 706 17 723 19
rect 706 13 709 17
rect 713 13 723 17
rect 1554 17 1560 19
rect 706 11 723 13
rect 4 -31 10 -29
rect 4 -35 5 -31
rect 9 -35 10 -31
rect 4 -37 10 -35
rect 14 -37 31 -29
rect 35 -31 52 -29
rect 35 -35 38 -31
rect 42 -35 52 -31
rect 35 -37 52 -35
rect 1554 13 1555 17
rect 1559 13 1560 17
rect 1554 11 1560 13
rect 1564 11 1581 19
rect 1585 17 1602 19
rect 1585 13 1588 17
rect 1592 13 1602 17
rect 2322 17 2328 19
rect 1585 11 1602 13
rect 602 -31 608 -29
rect 602 -35 603 -31
rect 607 -35 608 -31
rect 602 -37 608 -35
rect 612 -37 629 -29
rect 633 -31 650 -29
rect 633 -35 636 -31
rect 640 -35 650 -31
rect 633 -37 650 -35
rect 178 -51 184 -49
rect 178 -55 179 -51
rect 183 -55 184 -51
rect 178 -57 184 -55
rect 188 -57 205 -49
rect 209 -51 226 -49
rect 209 -55 212 -51
rect 216 -55 226 -51
rect 2322 13 2323 17
rect 2327 13 2328 17
rect 2322 11 2328 13
rect 2332 11 2349 19
rect 2353 17 2370 19
rect 2353 13 2356 17
rect 2360 13 2370 17
rect 2353 11 2370 13
rect 1481 -31 1487 -29
rect 1481 -35 1482 -31
rect 1486 -35 1487 -31
rect 1481 -37 1487 -35
rect 1491 -37 1508 -29
rect 1512 -31 1529 -29
rect 1512 -35 1515 -31
rect 1519 -35 1529 -31
rect 1512 -37 1529 -35
rect 776 -51 782 -49
rect 209 -57 226 -55
rect 776 -55 777 -51
rect 781 -55 782 -51
rect 776 -57 782 -55
rect 786 -57 803 -49
rect 807 -51 824 -49
rect 807 -55 810 -51
rect 814 -55 824 -51
rect 2249 -31 2255 -29
rect 2249 -35 2250 -31
rect 2254 -35 2255 -31
rect 2249 -37 2255 -35
rect 2259 -37 2276 -29
rect 2280 -31 2297 -29
rect 2280 -35 2283 -31
rect 2287 -35 2297 -31
rect 2280 -37 2297 -35
rect 1655 -51 1661 -49
rect 807 -57 824 -55
rect 1655 -55 1656 -51
rect 1660 -55 1661 -51
rect 1655 -57 1661 -55
rect 1665 -57 1682 -49
rect 1686 -51 1703 -49
rect 1686 -55 1689 -51
rect 1693 -55 1703 -51
rect 2423 -51 2429 -49
rect 1686 -57 1703 -55
rect 2423 -55 2424 -51
rect 2428 -55 2429 -51
rect 2423 -57 2429 -55
rect 2433 -57 2450 -49
rect 2454 -51 2471 -49
rect 2454 -55 2457 -51
rect 2461 -55 2471 -51
rect 2454 -57 2471 -55
rect 92 -92 98 -90
rect 92 -96 93 -92
rect 97 -96 98 -92
rect 92 -98 98 -96
rect 102 -98 119 -90
rect 123 -92 140 -90
rect 123 -96 126 -92
rect 130 -96 140 -92
rect 123 -98 140 -96
rect 690 -92 696 -90
rect 690 -96 691 -92
rect 695 -96 696 -92
rect 690 -98 696 -96
rect 700 -98 717 -90
rect 721 -92 738 -90
rect 721 -96 724 -92
rect 728 -96 738 -92
rect 721 -98 738 -96
rect 1569 -92 1575 -90
rect 1569 -96 1570 -92
rect 1574 -96 1575 -92
rect 1569 -98 1575 -96
rect 1579 -98 1596 -90
rect 1600 -92 1617 -90
rect 1600 -96 1603 -92
rect 1607 -96 1617 -92
rect 1600 -98 1617 -96
rect 2337 -92 2343 -90
rect 2337 -96 2338 -92
rect 2342 -96 2343 -92
rect 2337 -98 2343 -96
rect 2347 -98 2364 -90
rect 2368 -92 2385 -90
rect 2368 -96 2371 -92
rect 2375 -96 2385 -92
rect 2368 -98 2385 -96
rect 358 -286 364 -284
rect 358 -290 359 -286
rect 363 -290 364 -286
rect 358 -292 364 -290
rect 368 -292 385 -284
rect 389 -286 406 -284
rect 389 -290 392 -286
rect 396 -290 406 -286
rect 1101 -289 1107 -287
rect 389 -292 406 -290
rect 1101 -293 1102 -289
rect 1106 -293 1107 -289
rect 1101 -295 1107 -293
rect 1111 -295 1128 -287
rect 1132 -289 1149 -287
rect 1132 -293 1135 -289
rect 1139 -293 1149 -289
rect 1860 -289 1866 -287
rect 1132 -295 1149 -293
rect 48 -334 54 -332
rect 48 -338 49 -334
rect 53 -338 54 -334
rect 48 -340 54 -338
rect 58 -340 75 -332
rect 79 -334 96 -332
rect 79 -338 82 -334
rect 86 -338 96 -334
rect 79 -340 96 -338
rect 285 -334 291 -332
rect 285 -338 286 -334
rect 290 -338 291 -334
rect 285 -340 291 -338
rect 295 -340 312 -332
rect 316 -334 333 -332
rect 316 -338 319 -334
rect 323 -338 333 -334
rect 316 -340 333 -338
rect 1860 -293 1861 -289
rect 1865 -293 1866 -289
rect 1860 -295 1866 -293
rect 1870 -295 1887 -287
rect 1891 -289 1908 -287
rect 1891 -293 1894 -289
rect 1898 -293 1908 -289
rect 2596 -289 2602 -287
rect 1891 -295 1908 -293
rect 791 -337 797 -335
rect 791 -341 792 -337
rect 796 -341 797 -337
rect 791 -343 797 -341
rect 801 -343 818 -335
rect 822 -337 839 -335
rect 822 -341 825 -337
rect 829 -341 839 -337
rect 822 -343 839 -341
rect 1028 -337 1034 -335
rect 1028 -341 1029 -337
rect 1033 -341 1034 -337
rect 1028 -343 1034 -341
rect 1038 -343 1055 -335
rect 1059 -337 1076 -335
rect 1059 -341 1062 -337
rect 1066 -341 1076 -337
rect 1059 -343 1076 -341
rect 459 -354 465 -352
rect -25 -382 -19 -380
rect -25 -386 -24 -382
rect -20 -386 -19 -382
rect -25 -388 -19 -386
rect -15 -388 2 -380
rect 6 -382 23 -380
rect 6 -386 9 -382
rect 13 -386 23 -382
rect 6 -388 23 -386
rect 459 -358 460 -354
rect 464 -358 465 -354
rect 459 -360 465 -358
rect 469 -360 486 -352
rect 490 -354 507 -352
rect 490 -358 493 -354
rect 497 -358 507 -354
rect 490 -360 507 -358
rect 2596 -293 2597 -289
rect 2601 -293 2602 -289
rect 2596 -295 2602 -293
rect 2606 -295 2623 -287
rect 2627 -289 2644 -287
rect 2627 -293 2630 -289
rect 2634 -293 2644 -289
rect 2627 -295 2644 -293
rect 1550 -337 1556 -335
rect 1550 -341 1551 -337
rect 1555 -341 1556 -337
rect 1550 -343 1556 -341
rect 1560 -343 1577 -335
rect 1581 -337 1598 -335
rect 1581 -341 1584 -337
rect 1588 -341 1598 -337
rect 1581 -343 1598 -341
rect 1787 -337 1793 -335
rect 1787 -341 1788 -337
rect 1792 -341 1793 -337
rect 1787 -343 1793 -341
rect 1797 -343 1814 -335
rect 1818 -337 1835 -335
rect 1818 -341 1821 -337
rect 1825 -341 1835 -337
rect 1818 -343 1835 -341
rect 1202 -357 1208 -355
rect 718 -385 724 -383
rect 718 -389 719 -385
rect 723 -389 724 -385
rect 718 -391 724 -389
rect 728 -391 745 -383
rect 749 -385 766 -383
rect 749 -389 752 -385
rect 756 -389 766 -385
rect 749 -391 766 -389
rect 373 -395 379 -393
rect 373 -399 374 -395
rect 378 -399 379 -395
rect 149 -402 155 -400
rect 149 -406 150 -402
rect 154 -406 155 -402
rect 149 -408 155 -406
rect 159 -408 176 -400
rect 180 -402 197 -400
rect 373 -401 379 -399
rect 383 -401 400 -393
rect 404 -395 421 -393
rect 404 -399 407 -395
rect 411 -399 421 -395
rect 404 -401 421 -399
rect 180 -406 183 -402
rect 187 -406 197 -402
rect 180 -408 197 -406
rect 1202 -361 1203 -357
rect 1207 -361 1208 -357
rect 1202 -363 1208 -361
rect 1212 -363 1229 -355
rect 1233 -357 1250 -355
rect 1233 -361 1236 -357
rect 1240 -361 1250 -357
rect 1233 -363 1250 -361
rect 2286 -337 2292 -335
rect 2286 -341 2287 -337
rect 2291 -341 2292 -337
rect 2286 -343 2292 -341
rect 2296 -343 2313 -335
rect 2317 -337 2334 -335
rect 2317 -341 2320 -337
rect 2324 -341 2334 -337
rect 2317 -343 2334 -341
rect 2523 -337 2529 -335
rect 2523 -341 2524 -337
rect 2528 -341 2529 -337
rect 2523 -343 2529 -341
rect 2533 -343 2550 -335
rect 2554 -337 2571 -335
rect 2554 -341 2557 -337
rect 2561 -341 2571 -337
rect 2554 -343 2571 -341
rect 1961 -357 1967 -355
rect 1477 -385 1483 -383
rect 1477 -389 1478 -385
rect 1482 -389 1483 -385
rect 1477 -391 1483 -389
rect 1487 -391 1504 -383
rect 1508 -385 1525 -383
rect 1508 -389 1511 -385
rect 1515 -389 1525 -385
rect 1508 -391 1525 -389
rect 1116 -398 1122 -396
rect 1116 -402 1117 -398
rect 1121 -402 1122 -398
rect 892 -405 898 -403
rect 63 -443 69 -441
rect 63 -447 64 -443
rect 68 -447 69 -443
rect 63 -449 69 -447
rect 73 -449 90 -441
rect 94 -443 111 -441
rect 94 -447 97 -443
rect 101 -447 111 -443
rect 892 -409 893 -405
rect 897 -409 898 -405
rect 892 -411 898 -409
rect 902 -411 919 -403
rect 923 -405 940 -403
rect 1116 -404 1122 -402
rect 1126 -404 1143 -396
rect 1147 -398 1164 -396
rect 1147 -402 1150 -398
rect 1154 -402 1164 -398
rect 1147 -404 1164 -402
rect 923 -409 926 -405
rect 930 -409 940 -405
rect 923 -411 940 -409
rect 1961 -361 1962 -357
rect 1966 -361 1967 -357
rect 1961 -363 1967 -361
rect 1971 -363 1988 -355
rect 1992 -357 2009 -355
rect 1992 -361 1995 -357
rect 1999 -361 2009 -357
rect 1992 -363 2009 -361
rect 2697 -357 2703 -355
rect 2213 -385 2219 -383
rect 2213 -389 2214 -385
rect 2218 -389 2219 -385
rect 2213 -391 2219 -389
rect 2223 -391 2240 -383
rect 2244 -385 2261 -383
rect 2244 -389 2247 -385
rect 2251 -389 2261 -385
rect 2244 -391 2261 -389
rect 1875 -398 1881 -396
rect 1875 -402 1876 -398
rect 1880 -402 1881 -398
rect 1651 -405 1657 -403
rect 1651 -409 1652 -405
rect 1656 -409 1657 -405
rect 1651 -411 1657 -409
rect 1661 -411 1678 -403
rect 1682 -405 1699 -403
rect 1875 -404 1881 -402
rect 1885 -404 1902 -396
rect 1906 -398 1923 -396
rect 1906 -402 1909 -398
rect 1913 -402 1923 -398
rect 1906 -404 1923 -402
rect 1682 -409 1685 -405
rect 1689 -409 1699 -405
rect 1682 -411 1699 -409
rect 2697 -361 2698 -357
rect 2702 -361 2703 -357
rect 2697 -363 2703 -361
rect 2707 -363 2724 -355
rect 2728 -357 2745 -355
rect 2728 -361 2731 -357
rect 2735 -361 2745 -357
rect 2728 -363 2745 -361
rect 2611 -398 2617 -396
rect 2611 -402 2612 -398
rect 2616 -402 2617 -398
rect 2387 -405 2393 -403
rect 2387 -409 2388 -405
rect 2392 -409 2393 -405
rect 2387 -411 2393 -409
rect 2397 -411 2414 -403
rect 2418 -405 2435 -403
rect 2611 -404 2617 -402
rect 2621 -404 2638 -396
rect 2642 -398 2659 -396
rect 2642 -402 2645 -398
rect 2649 -402 2659 -398
rect 2642 -404 2659 -402
rect 2418 -409 2421 -405
rect 2425 -409 2435 -405
rect 2418 -411 2435 -409
rect 94 -449 111 -447
rect 806 -446 812 -444
rect 806 -450 807 -446
rect 811 -450 812 -446
rect 806 -452 812 -450
rect 816 -452 833 -444
rect 837 -446 854 -444
rect 837 -450 840 -446
rect 844 -450 854 -446
rect 837 -452 854 -450
rect 1565 -446 1571 -444
rect 1565 -450 1566 -446
rect 1570 -450 1571 -446
rect 1565 -452 1571 -450
rect 1575 -452 1592 -444
rect 1596 -446 1613 -444
rect 1596 -450 1599 -446
rect 1603 -450 1613 -446
rect 1596 -452 1613 -450
rect 2301 -446 2307 -444
rect 2301 -450 2302 -446
rect 2306 -450 2307 -446
rect 2301 -452 2307 -450
rect 2311 -452 2328 -444
rect 2332 -446 2349 -444
rect 2332 -450 2335 -446
rect 2339 -450 2349 -446
rect 2332 -452 2349 -450
rect 345 -501 351 -499
rect 345 -505 346 -501
rect 350 -505 351 -501
rect 345 -507 351 -505
rect 355 -507 372 -499
rect 376 -501 393 -499
rect 376 -505 379 -501
rect 383 -505 393 -501
rect 376 -507 393 -505
rect 411 -501 417 -499
rect 411 -505 412 -501
rect 416 -505 417 -501
rect 411 -507 417 -505
rect 421 -501 427 -499
rect 421 -505 422 -501
rect 426 -505 427 -501
rect 421 -507 427 -505
rect 504 -504 510 -502
rect 504 -508 505 -504
rect 509 -508 510 -504
rect 504 -510 510 -508
rect 514 -504 531 -502
rect 514 -508 515 -504
rect 519 -508 531 -504
rect 514 -510 531 -508
rect 535 -504 552 -502
rect 535 -508 538 -504
rect 542 -508 552 -504
rect 535 -510 552 -508
rect 572 -504 578 -502
rect 572 -508 573 -504
rect 577 -508 578 -504
rect 572 -510 578 -508
rect 582 -504 588 -502
rect 582 -508 583 -504
rect 587 -508 588 -504
rect 1088 -504 1094 -502
rect 1088 -508 1089 -504
rect 1093 -508 1094 -504
rect 582 -510 588 -508
rect 1088 -510 1094 -508
rect 1098 -510 1115 -502
rect 1119 -504 1136 -502
rect 1119 -508 1122 -504
rect 1126 -508 1136 -504
rect 1119 -510 1136 -508
rect 1154 -504 1160 -502
rect 1154 -508 1155 -504
rect 1159 -508 1160 -504
rect 1154 -510 1160 -508
rect 1164 -504 1170 -502
rect 1164 -508 1165 -504
rect 1169 -508 1170 -504
rect 1847 -504 1853 -502
rect 1164 -510 1170 -508
rect 1247 -507 1253 -505
rect 1247 -511 1248 -507
rect 1252 -511 1253 -507
rect 1247 -513 1253 -511
rect 1257 -507 1274 -505
rect 1257 -511 1258 -507
rect 1262 -511 1274 -507
rect 1257 -513 1274 -511
rect 1278 -507 1295 -505
rect 1278 -511 1281 -507
rect 1285 -511 1295 -507
rect 1278 -513 1295 -511
rect 1315 -507 1321 -505
rect 1315 -511 1316 -507
rect 1320 -511 1321 -507
rect 1315 -513 1321 -511
rect 1325 -507 1331 -505
rect 1325 -511 1326 -507
rect 1330 -511 1331 -507
rect 1847 -508 1848 -504
rect 1852 -508 1853 -504
rect 1325 -513 1331 -511
rect 1847 -510 1853 -508
rect 1857 -510 1874 -502
rect 1878 -504 1895 -502
rect 1878 -508 1881 -504
rect 1885 -508 1895 -504
rect 1878 -510 1895 -508
rect 1913 -504 1919 -502
rect 1913 -508 1914 -504
rect 1918 -508 1919 -504
rect 1913 -510 1919 -508
rect 1923 -504 1929 -502
rect 1923 -508 1924 -504
rect 1928 -508 1929 -504
rect 2583 -504 2589 -502
rect 1923 -510 1929 -508
rect 2006 -507 2012 -505
rect 2006 -511 2007 -507
rect 2011 -511 2012 -507
rect 2006 -513 2012 -511
rect 2016 -507 2033 -505
rect 2016 -511 2017 -507
rect 2021 -511 2033 -507
rect 2016 -513 2033 -511
rect 2037 -507 2054 -505
rect 2037 -511 2040 -507
rect 2044 -511 2054 -507
rect 2037 -513 2054 -511
rect 2074 -507 2080 -505
rect 2074 -511 2075 -507
rect 2079 -511 2080 -507
rect 2074 -513 2080 -511
rect 2084 -507 2090 -505
rect 2084 -511 2085 -507
rect 2089 -511 2090 -507
rect 2583 -508 2584 -504
rect 2588 -508 2589 -504
rect 2084 -513 2090 -511
rect 2583 -510 2589 -508
rect 2593 -510 2610 -502
rect 2614 -504 2631 -502
rect 2614 -508 2617 -504
rect 2621 -508 2631 -504
rect 2614 -510 2631 -508
rect 2649 -504 2655 -502
rect 2649 -508 2650 -504
rect 2654 -508 2655 -504
rect 2649 -510 2655 -508
rect 2659 -504 2665 -502
rect 2659 -508 2660 -504
rect 2664 -508 2665 -504
rect 2659 -510 2665 -508
rect 2742 -507 2748 -505
rect 2742 -511 2743 -507
rect 2747 -511 2748 -507
rect 2742 -513 2748 -511
rect 2752 -507 2769 -505
rect 2752 -511 2753 -507
rect 2757 -511 2769 -507
rect 2752 -513 2769 -511
rect 2773 -507 2790 -505
rect 2773 -511 2776 -507
rect 2780 -511 2790 -507
rect 2773 -513 2790 -511
rect 2810 -507 2816 -505
rect 2810 -511 2811 -507
rect 2815 -511 2816 -507
rect 2810 -513 2816 -511
rect 2820 -507 2826 -505
rect 2820 -511 2821 -507
rect 2825 -511 2826 -507
rect 2820 -513 2826 -511
rect 34 -552 40 -550
rect 34 -556 35 -552
rect 39 -556 40 -552
rect 34 -558 40 -556
rect 44 -558 61 -550
rect 65 -552 82 -550
rect 65 -556 68 -552
rect 72 -556 82 -552
rect 65 -558 82 -556
rect 100 -552 106 -550
rect 100 -556 101 -552
rect 105 -556 106 -552
rect 100 -558 106 -556
rect 110 -552 116 -550
rect 110 -556 111 -552
rect 115 -556 116 -552
rect 110 -558 116 -556
rect 777 -555 783 -553
rect 777 -559 778 -555
rect 782 -559 783 -555
rect 777 -561 783 -559
rect 787 -561 804 -553
rect 808 -555 825 -553
rect 808 -559 811 -555
rect 815 -559 825 -555
rect 808 -561 825 -559
rect 843 -555 849 -553
rect 843 -559 844 -555
rect 848 -559 849 -555
rect 843 -561 849 -559
rect 853 -555 859 -553
rect 853 -559 854 -555
rect 858 -559 859 -555
rect 853 -561 859 -559
rect 1536 -555 1542 -553
rect 1536 -559 1537 -555
rect 1541 -559 1542 -555
rect 1536 -561 1542 -559
rect 1546 -561 1563 -553
rect 1567 -555 1584 -553
rect 1567 -559 1570 -555
rect 1574 -559 1584 -555
rect 1567 -561 1584 -559
rect 1602 -555 1608 -553
rect 1602 -559 1603 -555
rect 1607 -559 1608 -555
rect 1602 -561 1608 -559
rect 1612 -555 1618 -553
rect 1612 -559 1613 -555
rect 1617 -559 1618 -555
rect 1612 -561 1618 -559
rect 2272 -555 2278 -553
rect 2272 -559 2273 -555
rect 2277 -559 2278 -555
rect 2272 -561 2278 -559
rect 2282 -561 2299 -553
rect 2303 -555 2320 -553
rect 2303 -559 2306 -555
rect 2310 -559 2320 -555
rect 2303 -561 2320 -559
rect 2338 -555 2344 -553
rect 2338 -559 2339 -555
rect 2343 -559 2344 -555
rect 2338 -561 2344 -559
rect 2348 -555 2354 -553
rect 2348 -559 2349 -555
rect 2353 -559 2354 -555
rect 2348 -561 2354 -559
<< pdiffusion >>
rect 77 62 83 64
rect 77 58 78 62
rect 82 58 83 62
rect 77 56 83 58
rect 87 62 104 64
rect 87 58 88 62
rect 92 58 104 62
rect 87 56 104 58
rect 108 62 125 64
rect 108 58 111 62
rect 115 58 125 62
rect 108 56 125 58
rect 675 62 681 64
rect 675 58 676 62
rect 680 58 681 62
rect 675 56 681 58
rect 685 62 702 64
rect 685 58 686 62
rect 690 58 702 62
rect 685 56 702 58
rect 706 62 723 64
rect 706 58 709 62
rect 713 58 723 62
rect 706 56 723 58
rect 1554 62 1560 64
rect 1554 58 1555 62
rect 1559 58 1560 62
rect 1554 56 1560 58
rect 1564 62 1581 64
rect 1564 58 1565 62
rect 1569 58 1581 62
rect 1564 56 1581 58
rect 1585 62 1602 64
rect 1585 58 1588 62
rect 1592 58 1602 62
rect 1585 56 1602 58
rect 2322 62 2328 64
rect 2322 58 2323 62
rect 2327 58 2328 62
rect 2322 56 2328 58
rect 2332 62 2349 64
rect 2332 58 2333 62
rect 2337 58 2349 62
rect 2332 56 2349 58
rect 2353 62 2370 64
rect 2353 58 2356 62
rect 2360 58 2370 62
rect 2353 56 2370 58
rect 4 14 10 16
rect 4 10 5 14
rect 9 10 10 14
rect 4 8 10 10
rect 14 14 31 16
rect 14 10 15 14
rect 19 10 31 14
rect 14 8 31 10
rect 35 14 52 16
rect 35 10 38 14
rect 42 10 52 14
rect 602 14 608 16
rect 35 8 52 10
rect 602 10 603 14
rect 607 10 608 14
rect 602 8 608 10
rect 612 14 629 16
rect 612 10 613 14
rect 617 10 629 14
rect 612 8 629 10
rect 633 14 650 16
rect 633 10 636 14
rect 640 10 650 14
rect 1481 14 1487 16
rect 633 8 650 10
rect 178 -6 184 -4
rect 178 -10 179 -6
rect 183 -10 184 -6
rect 178 -12 184 -10
rect 188 -6 205 -4
rect 188 -10 189 -6
rect 193 -10 205 -6
rect 188 -12 205 -10
rect 209 -6 226 -4
rect 209 -10 212 -6
rect 216 -10 226 -6
rect 209 -12 226 -10
rect 92 -47 98 -45
rect 92 -51 93 -47
rect 97 -51 98 -47
rect 92 -53 98 -51
rect 102 -47 119 -45
rect 102 -51 103 -47
rect 107 -51 119 -47
rect 102 -53 119 -51
rect 123 -47 140 -45
rect 123 -51 126 -47
rect 130 -51 140 -47
rect 1481 10 1482 14
rect 1486 10 1487 14
rect 1481 8 1487 10
rect 1491 14 1508 16
rect 1491 10 1492 14
rect 1496 10 1508 14
rect 1491 8 1508 10
rect 1512 14 1529 16
rect 1512 10 1515 14
rect 1519 10 1529 14
rect 2249 14 2255 16
rect 1512 8 1529 10
rect 776 -6 782 -4
rect 776 -10 777 -6
rect 781 -10 782 -6
rect 776 -12 782 -10
rect 786 -6 803 -4
rect 786 -10 787 -6
rect 791 -10 803 -6
rect 786 -12 803 -10
rect 807 -6 824 -4
rect 807 -10 810 -6
rect 814 -10 824 -6
rect 807 -12 824 -10
rect 690 -47 696 -45
rect 123 -53 140 -51
rect 690 -51 691 -47
rect 695 -51 696 -47
rect 690 -53 696 -51
rect 700 -47 717 -45
rect 700 -51 701 -47
rect 705 -51 717 -47
rect 700 -53 717 -51
rect 721 -47 738 -45
rect 721 -51 724 -47
rect 728 -51 738 -47
rect 2249 10 2250 14
rect 2254 10 2255 14
rect 2249 8 2255 10
rect 2259 14 2276 16
rect 2259 10 2260 14
rect 2264 10 2276 14
rect 2259 8 2276 10
rect 2280 14 2297 16
rect 2280 10 2283 14
rect 2287 10 2297 14
rect 2280 8 2297 10
rect 1655 -6 1661 -4
rect 1655 -10 1656 -6
rect 1660 -10 1661 -6
rect 1655 -12 1661 -10
rect 1665 -6 1682 -4
rect 1665 -10 1666 -6
rect 1670 -10 1682 -6
rect 1665 -12 1682 -10
rect 1686 -6 1703 -4
rect 1686 -10 1689 -6
rect 1693 -10 1703 -6
rect 1686 -12 1703 -10
rect 1569 -47 1575 -45
rect 721 -53 738 -51
rect 1569 -51 1570 -47
rect 1574 -51 1575 -47
rect 1569 -53 1575 -51
rect 1579 -47 1596 -45
rect 1579 -51 1580 -47
rect 1584 -51 1596 -47
rect 1579 -53 1596 -51
rect 1600 -47 1617 -45
rect 1600 -51 1603 -47
rect 1607 -51 1617 -47
rect 2423 -6 2429 -4
rect 2423 -10 2424 -6
rect 2428 -10 2429 -6
rect 2423 -12 2429 -10
rect 2433 -6 2450 -4
rect 2433 -10 2434 -6
rect 2438 -10 2450 -6
rect 2433 -12 2450 -10
rect 2454 -6 2471 -4
rect 2454 -10 2457 -6
rect 2461 -10 2471 -6
rect 2454 -12 2471 -10
rect 2337 -47 2343 -45
rect 1600 -53 1617 -51
rect 2337 -51 2338 -47
rect 2342 -51 2343 -47
rect 2337 -53 2343 -51
rect 2347 -47 2364 -45
rect 2347 -51 2348 -47
rect 2352 -51 2364 -47
rect 2347 -53 2364 -51
rect 2368 -47 2385 -45
rect 2368 -51 2371 -47
rect 2375 -51 2385 -47
rect 2368 -53 2385 -51
rect 358 -241 364 -239
rect 358 -245 359 -241
rect 363 -245 364 -241
rect 358 -247 364 -245
rect 368 -241 385 -239
rect 368 -245 369 -241
rect 373 -245 385 -241
rect 368 -247 385 -245
rect 389 -241 406 -239
rect 389 -245 392 -241
rect 396 -245 406 -241
rect 389 -247 406 -245
rect 1101 -244 1107 -242
rect 1101 -248 1102 -244
rect 1106 -248 1107 -244
rect 1101 -250 1107 -248
rect 1111 -244 1128 -242
rect 1111 -248 1112 -244
rect 1116 -248 1128 -244
rect 1111 -250 1128 -248
rect 1132 -244 1149 -242
rect 1132 -248 1135 -244
rect 1139 -248 1149 -244
rect 1132 -250 1149 -248
rect 1860 -244 1866 -242
rect 1860 -248 1861 -244
rect 1865 -248 1866 -244
rect 1860 -250 1866 -248
rect 1870 -244 1887 -242
rect 1870 -248 1871 -244
rect 1875 -248 1887 -244
rect 1870 -250 1887 -248
rect 1891 -244 1908 -242
rect 1891 -248 1894 -244
rect 1898 -248 1908 -244
rect 1891 -250 1908 -248
rect 2596 -244 2602 -242
rect 2596 -248 2597 -244
rect 2601 -248 2602 -244
rect 2596 -250 2602 -248
rect 2606 -244 2623 -242
rect 2606 -248 2607 -244
rect 2611 -248 2623 -244
rect 2606 -250 2623 -248
rect 2627 -244 2644 -242
rect 2627 -248 2630 -244
rect 2634 -248 2644 -244
rect 2627 -250 2644 -248
rect 48 -289 54 -287
rect 48 -293 49 -289
rect 53 -293 54 -289
rect 48 -295 54 -293
rect 58 -289 75 -287
rect 58 -293 59 -289
rect 63 -293 75 -289
rect 58 -295 75 -293
rect 79 -289 96 -287
rect 79 -293 82 -289
rect 86 -293 96 -289
rect 79 -295 96 -293
rect 285 -289 291 -287
rect 285 -293 286 -289
rect 290 -293 291 -289
rect 285 -295 291 -293
rect 295 -289 312 -287
rect 295 -293 296 -289
rect 300 -293 312 -289
rect 295 -295 312 -293
rect 316 -289 333 -287
rect 316 -293 319 -289
rect 323 -293 333 -289
rect 791 -292 797 -290
rect 316 -295 333 -293
rect 791 -296 792 -292
rect 796 -296 797 -292
rect 791 -298 797 -296
rect 801 -292 818 -290
rect 801 -296 802 -292
rect 806 -296 818 -292
rect 801 -298 818 -296
rect 822 -292 839 -290
rect 822 -296 825 -292
rect 829 -296 839 -292
rect 822 -298 839 -296
rect 1028 -292 1034 -290
rect 1028 -296 1029 -292
rect 1033 -296 1034 -292
rect 1028 -298 1034 -296
rect 1038 -292 1055 -290
rect 1038 -296 1039 -292
rect 1043 -296 1055 -292
rect 1038 -298 1055 -296
rect 1059 -292 1076 -290
rect 1059 -296 1062 -292
rect 1066 -296 1076 -292
rect 1550 -292 1556 -290
rect 1059 -298 1076 -296
rect 459 -309 465 -307
rect 459 -313 460 -309
rect 464 -313 465 -309
rect 459 -315 465 -313
rect 469 -309 486 -307
rect 469 -313 470 -309
rect 474 -313 486 -309
rect 469 -315 486 -313
rect 490 -309 507 -307
rect 490 -313 493 -309
rect 497 -313 507 -309
rect 490 -315 507 -313
rect -25 -337 -19 -335
rect -25 -341 -24 -337
rect -20 -341 -19 -337
rect -25 -343 -19 -341
rect -15 -337 2 -335
rect -15 -341 -14 -337
rect -10 -341 2 -337
rect -15 -343 2 -341
rect 6 -337 23 -335
rect 6 -341 9 -337
rect 13 -341 23 -337
rect 6 -343 23 -341
rect 373 -350 379 -348
rect 373 -354 374 -350
rect 378 -354 379 -350
rect 149 -357 155 -355
rect 149 -361 150 -357
rect 154 -361 155 -357
rect 149 -363 155 -361
rect 159 -357 176 -355
rect 159 -361 160 -357
rect 164 -361 176 -357
rect 159 -363 176 -361
rect 180 -357 197 -355
rect 373 -356 379 -354
rect 383 -350 400 -348
rect 383 -354 384 -350
rect 388 -354 400 -350
rect 383 -356 400 -354
rect 404 -350 421 -348
rect 404 -354 407 -350
rect 411 -354 421 -350
rect 1550 -296 1551 -292
rect 1555 -296 1556 -292
rect 1550 -298 1556 -296
rect 1560 -292 1577 -290
rect 1560 -296 1561 -292
rect 1565 -296 1577 -292
rect 1560 -298 1577 -296
rect 1581 -292 1598 -290
rect 1581 -296 1584 -292
rect 1588 -296 1598 -292
rect 1581 -298 1598 -296
rect 1787 -292 1793 -290
rect 1787 -296 1788 -292
rect 1792 -296 1793 -292
rect 1787 -298 1793 -296
rect 1797 -292 1814 -290
rect 1797 -296 1798 -292
rect 1802 -296 1814 -292
rect 1797 -298 1814 -296
rect 1818 -292 1835 -290
rect 1818 -296 1821 -292
rect 1825 -296 1835 -292
rect 2286 -292 2292 -290
rect 1818 -298 1835 -296
rect 1202 -312 1208 -310
rect 1202 -316 1203 -312
rect 1207 -316 1208 -312
rect 1202 -318 1208 -316
rect 1212 -312 1229 -310
rect 1212 -316 1213 -312
rect 1217 -316 1229 -312
rect 1212 -318 1229 -316
rect 1233 -312 1250 -310
rect 1233 -316 1236 -312
rect 1240 -316 1250 -312
rect 1233 -318 1250 -316
rect 718 -340 724 -338
rect 718 -344 719 -340
rect 723 -344 724 -340
rect 718 -346 724 -344
rect 728 -340 745 -338
rect 728 -344 729 -340
rect 733 -344 745 -340
rect 728 -346 745 -344
rect 749 -340 766 -338
rect 749 -344 752 -340
rect 756 -344 766 -340
rect 749 -346 766 -344
rect 404 -356 421 -354
rect 180 -361 183 -357
rect 187 -361 197 -357
rect 180 -363 197 -361
rect 63 -398 69 -396
rect 63 -402 64 -398
rect 68 -402 69 -398
rect 63 -404 69 -402
rect 73 -398 90 -396
rect 73 -402 74 -398
rect 78 -402 90 -398
rect 73 -404 90 -402
rect 94 -398 111 -396
rect 94 -402 97 -398
rect 101 -402 111 -398
rect 1116 -353 1122 -351
rect 1116 -357 1117 -353
rect 1121 -357 1122 -353
rect 892 -360 898 -358
rect 892 -364 893 -360
rect 897 -364 898 -360
rect 892 -366 898 -364
rect 902 -360 919 -358
rect 902 -364 903 -360
rect 907 -364 919 -360
rect 902 -366 919 -364
rect 923 -360 940 -358
rect 1116 -359 1122 -357
rect 1126 -353 1143 -351
rect 1126 -357 1127 -353
rect 1131 -357 1143 -353
rect 1126 -359 1143 -357
rect 1147 -353 1164 -351
rect 1147 -357 1150 -353
rect 1154 -357 1164 -353
rect 2286 -296 2287 -292
rect 2291 -296 2292 -292
rect 2286 -298 2292 -296
rect 2296 -292 2313 -290
rect 2296 -296 2297 -292
rect 2301 -296 2313 -292
rect 2296 -298 2313 -296
rect 2317 -292 2334 -290
rect 2317 -296 2320 -292
rect 2324 -296 2334 -292
rect 2317 -298 2334 -296
rect 2523 -292 2529 -290
rect 2523 -296 2524 -292
rect 2528 -296 2529 -292
rect 2523 -298 2529 -296
rect 2533 -292 2550 -290
rect 2533 -296 2534 -292
rect 2538 -296 2550 -292
rect 2533 -298 2550 -296
rect 2554 -292 2571 -290
rect 2554 -296 2557 -292
rect 2561 -296 2571 -292
rect 2554 -298 2571 -296
rect 1961 -312 1967 -310
rect 1961 -316 1962 -312
rect 1966 -316 1967 -312
rect 1961 -318 1967 -316
rect 1971 -312 1988 -310
rect 1971 -316 1972 -312
rect 1976 -316 1988 -312
rect 1971 -318 1988 -316
rect 1992 -312 2009 -310
rect 1992 -316 1995 -312
rect 1999 -316 2009 -312
rect 1992 -318 2009 -316
rect 1477 -340 1483 -338
rect 1477 -344 1478 -340
rect 1482 -344 1483 -340
rect 1477 -346 1483 -344
rect 1487 -340 1504 -338
rect 1487 -344 1488 -340
rect 1492 -344 1504 -340
rect 1487 -346 1504 -344
rect 1508 -340 1525 -338
rect 1508 -344 1511 -340
rect 1515 -344 1525 -340
rect 1508 -346 1525 -344
rect 1147 -359 1164 -357
rect 923 -364 926 -360
rect 930 -364 940 -360
rect 923 -366 940 -364
rect 94 -404 111 -402
rect 806 -401 812 -399
rect 806 -405 807 -401
rect 811 -405 812 -401
rect 806 -407 812 -405
rect 816 -401 833 -399
rect 816 -405 817 -401
rect 821 -405 833 -401
rect 816 -407 833 -405
rect 837 -401 854 -399
rect 837 -405 840 -401
rect 844 -405 854 -401
rect 1875 -353 1881 -351
rect 1875 -357 1876 -353
rect 1880 -357 1881 -353
rect 1651 -360 1657 -358
rect 1651 -364 1652 -360
rect 1656 -364 1657 -360
rect 1651 -366 1657 -364
rect 1661 -360 1678 -358
rect 1661 -364 1662 -360
rect 1666 -364 1678 -360
rect 1661 -366 1678 -364
rect 1682 -360 1699 -358
rect 1875 -359 1881 -357
rect 1885 -353 1902 -351
rect 1885 -357 1886 -353
rect 1890 -357 1902 -353
rect 1885 -359 1902 -357
rect 1906 -353 1923 -351
rect 1906 -357 1909 -353
rect 1913 -357 1923 -353
rect 2697 -312 2703 -310
rect 2697 -316 2698 -312
rect 2702 -316 2703 -312
rect 2697 -318 2703 -316
rect 2707 -312 2724 -310
rect 2707 -316 2708 -312
rect 2712 -316 2724 -312
rect 2707 -318 2724 -316
rect 2728 -312 2745 -310
rect 2728 -316 2731 -312
rect 2735 -316 2745 -312
rect 2728 -318 2745 -316
rect 2213 -340 2219 -338
rect 2213 -344 2214 -340
rect 2218 -344 2219 -340
rect 2213 -346 2219 -344
rect 2223 -340 2240 -338
rect 2223 -344 2224 -340
rect 2228 -344 2240 -340
rect 2223 -346 2240 -344
rect 2244 -340 2261 -338
rect 2244 -344 2247 -340
rect 2251 -344 2261 -340
rect 2244 -346 2261 -344
rect 1906 -359 1923 -357
rect 1682 -364 1685 -360
rect 1689 -364 1699 -360
rect 1682 -366 1699 -364
rect 837 -407 854 -405
rect 1565 -401 1571 -399
rect 1565 -405 1566 -401
rect 1570 -405 1571 -401
rect 1565 -407 1571 -405
rect 1575 -401 1592 -399
rect 1575 -405 1576 -401
rect 1580 -405 1592 -401
rect 1575 -407 1592 -405
rect 1596 -401 1613 -399
rect 1596 -405 1599 -401
rect 1603 -405 1613 -401
rect 2611 -353 2617 -351
rect 2611 -357 2612 -353
rect 2616 -357 2617 -353
rect 2387 -360 2393 -358
rect 2387 -364 2388 -360
rect 2392 -364 2393 -360
rect 2387 -366 2393 -364
rect 2397 -360 2414 -358
rect 2397 -364 2398 -360
rect 2402 -364 2414 -360
rect 2397 -366 2414 -364
rect 2418 -360 2435 -358
rect 2611 -359 2617 -357
rect 2621 -353 2638 -351
rect 2621 -357 2622 -353
rect 2626 -357 2638 -353
rect 2621 -359 2638 -357
rect 2642 -353 2659 -351
rect 2642 -357 2645 -353
rect 2649 -357 2659 -353
rect 2642 -359 2659 -357
rect 2418 -364 2421 -360
rect 2425 -364 2435 -360
rect 2418 -366 2435 -364
rect 1596 -407 1613 -405
rect 2301 -401 2307 -399
rect 2301 -405 2302 -401
rect 2306 -405 2307 -401
rect 2301 -407 2307 -405
rect 2311 -401 2328 -399
rect 2311 -405 2312 -401
rect 2316 -405 2328 -401
rect 2311 -407 2328 -405
rect 2332 -401 2349 -399
rect 2332 -405 2335 -401
rect 2339 -405 2349 -401
rect 2332 -407 2349 -405
rect 345 -456 351 -454
rect 345 -460 346 -456
rect 350 -460 351 -456
rect 345 -462 351 -460
rect 355 -456 372 -454
rect 355 -460 356 -456
rect 360 -460 372 -456
rect 355 -462 372 -460
rect 376 -456 393 -454
rect 376 -460 379 -456
rect 383 -460 393 -456
rect 376 -462 393 -460
rect 411 -456 417 -454
rect 411 -460 412 -456
rect 416 -460 417 -456
rect 411 -462 417 -460
rect 421 -456 427 -454
rect 421 -460 422 -456
rect 426 -460 427 -456
rect 421 -462 427 -460
rect 504 -456 510 -454
rect 504 -460 505 -456
rect 509 -460 510 -456
rect 504 -462 510 -460
rect 514 -462 531 -454
rect 535 -456 552 -454
rect 535 -460 540 -456
rect 544 -460 552 -456
rect 535 -462 552 -460
rect 572 -456 578 -454
rect 572 -460 573 -456
rect 577 -460 578 -456
rect 572 -462 578 -460
rect 582 -456 588 -454
rect 582 -460 583 -456
rect 587 -460 588 -456
rect 1088 -459 1094 -457
rect 582 -462 588 -460
rect 34 -507 40 -505
rect 34 -511 35 -507
rect 39 -511 40 -507
rect 34 -513 40 -511
rect 44 -507 61 -505
rect 44 -511 45 -507
rect 49 -511 61 -507
rect 44 -513 61 -511
rect 65 -507 82 -505
rect 65 -511 68 -507
rect 72 -511 82 -507
rect 65 -513 82 -511
rect 100 -507 106 -505
rect 100 -511 101 -507
rect 105 -511 106 -507
rect 100 -513 106 -511
rect 110 -507 116 -505
rect 1088 -463 1089 -459
rect 1093 -463 1094 -459
rect 1088 -465 1094 -463
rect 1098 -459 1115 -457
rect 1098 -463 1099 -459
rect 1103 -463 1115 -459
rect 1098 -465 1115 -463
rect 1119 -459 1136 -457
rect 1119 -463 1122 -459
rect 1126 -463 1136 -459
rect 1119 -465 1136 -463
rect 1154 -459 1160 -457
rect 1154 -463 1155 -459
rect 1159 -463 1160 -459
rect 1154 -465 1160 -463
rect 1164 -459 1170 -457
rect 1164 -463 1165 -459
rect 1169 -463 1170 -459
rect 1164 -465 1170 -463
rect 1247 -459 1253 -457
rect 1247 -463 1248 -459
rect 1252 -463 1253 -459
rect 1247 -465 1253 -463
rect 1257 -465 1274 -457
rect 1278 -459 1295 -457
rect 1278 -463 1283 -459
rect 1287 -463 1295 -459
rect 1278 -465 1295 -463
rect 1315 -459 1321 -457
rect 1315 -463 1316 -459
rect 1320 -463 1321 -459
rect 1315 -465 1321 -463
rect 1325 -459 1331 -457
rect 1325 -463 1326 -459
rect 1330 -463 1331 -459
rect 1847 -459 1853 -457
rect 1325 -465 1331 -463
rect 1847 -463 1848 -459
rect 1852 -463 1853 -459
rect 1847 -465 1853 -463
rect 1857 -459 1874 -457
rect 1857 -463 1858 -459
rect 1862 -463 1874 -459
rect 1857 -465 1874 -463
rect 1878 -459 1895 -457
rect 1878 -463 1881 -459
rect 1885 -463 1895 -459
rect 1878 -465 1895 -463
rect 1913 -459 1919 -457
rect 1913 -463 1914 -459
rect 1918 -463 1919 -459
rect 1913 -465 1919 -463
rect 1923 -459 1929 -457
rect 1923 -463 1924 -459
rect 1928 -463 1929 -459
rect 1923 -465 1929 -463
rect 2006 -459 2012 -457
rect 2006 -463 2007 -459
rect 2011 -463 2012 -459
rect 2006 -465 2012 -463
rect 2016 -465 2033 -457
rect 2037 -459 2054 -457
rect 2037 -463 2042 -459
rect 2046 -463 2054 -459
rect 2037 -465 2054 -463
rect 2074 -459 2080 -457
rect 2074 -463 2075 -459
rect 2079 -463 2080 -459
rect 2074 -465 2080 -463
rect 2084 -459 2090 -457
rect 2084 -463 2085 -459
rect 2089 -463 2090 -459
rect 2583 -459 2589 -457
rect 2084 -465 2090 -463
rect 2583 -463 2584 -459
rect 2588 -463 2589 -459
rect 2583 -465 2589 -463
rect 2593 -459 2610 -457
rect 2593 -463 2594 -459
rect 2598 -463 2610 -459
rect 2593 -465 2610 -463
rect 2614 -459 2631 -457
rect 2614 -463 2617 -459
rect 2621 -463 2631 -459
rect 2614 -465 2631 -463
rect 2649 -459 2655 -457
rect 2649 -463 2650 -459
rect 2654 -463 2655 -459
rect 2649 -465 2655 -463
rect 2659 -459 2665 -457
rect 2659 -463 2660 -459
rect 2664 -463 2665 -459
rect 2659 -465 2665 -463
rect 2742 -459 2748 -457
rect 2742 -463 2743 -459
rect 2747 -463 2748 -459
rect 2742 -465 2748 -463
rect 2752 -465 2769 -457
rect 2773 -459 2790 -457
rect 2773 -463 2778 -459
rect 2782 -463 2790 -459
rect 2773 -465 2790 -463
rect 2810 -459 2816 -457
rect 2810 -463 2811 -459
rect 2815 -463 2816 -459
rect 2810 -465 2816 -463
rect 2820 -459 2826 -457
rect 2820 -463 2821 -459
rect 2825 -463 2826 -459
rect 2820 -465 2826 -463
rect 110 -511 111 -507
rect 115 -511 116 -507
rect 777 -510 783 -508
rect 110 -513 116 -511
rect 777 -514 778 -510
rect 782 -514 783 -510
rect 777 -516 783 -514
rect 787 -510 804 -508
rect 787 -514 788 -510
rect 792 -514 804 -510
rect 787 -516 804 -514
rect 808 -510 825 -508
rect 808 -514 811 -510
rect 815 -514 825 -510
rect 808 -516 825 -514
rect 843 -510 849 -508
rect 843 -514 844 -510
rect 848 -514 849 -510
rect 843 -516 849 -514
rect 853 -510 859 -508
rect 853 -514 854 -510
rect 858 -514 859 -510
rect 1536 -510 1542 -508
rect 853 -516 859 -514
rect 1536 -514 1537 -510
rect 1541 -514 1542 -510
rect 1536 -516 1542 -514
rect 1546 -510 1563 -508
rect 1546 -514 1547 -510
rect 1551 -514 1563 -510
rect 1546 -516 1563 -514
rect 1567 -510 1584 -508
rect 1567 -514 1570 -510
rect 1574 -514 1584 -510
rect 1567 -516 1584 -514
rect 1602 -510 1608 -508
rect 1602 -514 1603 -510
rect 1607 -514 1608 -510
rect 1602 -516 1608 -514
rect 1612 -510 1618 -508
rect 1612 -514 1613 -510
rect 1617 -514 1618 -510
rect 2272 -510 2278 -508
rect 1612 -516 1618 -514
rect 2272 -514 2273 -510
rect 2277 -514 2278 -510
rect 2272 -516 2278 -514
rect 2282 -510 2299 -508
rect 2282 -514 2283 -510
rect 2287 -514 2299 -510
rect 2282 -516 2299 -514
rect 2303 -510 2320 -508
rect 2303 -514 2306 -510
rect 2310 -514 2320 -510
rect 2303 -516 2320 -514
rect 2338 -510 2344 -508
rect 2338 -514 2339 -510
rect 2343 -514 2344 -510
rect 2338 -516 2344 -514
rect 2348 -510 2354 -508
rect 2348 -514 2349 -510
rect 2353 -514 2354 -510
rect 2348 -516 2354 -514
<< ndcontact >>
rect 78 13 82 17
rect 111 13 115 17
rect 676 13 680 17
rect 709 13 713 17
rect 5 -35 9 -31
rect 38 -35 42 -31
rect 1555 13 1559 17
rect 1588 13 1592 17
rect 603 -35 607 -31
rect 636 -35 640 -31
rect 179 -55 183 -51
rect 212 -55 216 -51
rect 2323 13 2327 17
rect 2356 13 2360 17
rect 1482 -35 1486 -31
rect 1515 -35 1519 -31
rect 777 -55 781 -51
rect 810 -55 814 -51
rect 2250 -35 2254 -31
rect 2283 -35 2287 -31
rect 1656 -55 1660 -51
rect 1689 -55 1693 -51
rect 2424 -55 2428 -51
rect 2457 -55 2461 -51
rect 93 -96 97 -92
rect 126 -96 130 -92
rect 691 -96 695 -92
rect 724 -96 728 -92
rect 1570 -96 1574 -92
rect 1603 -96 1607 -92
rect 2338 -96 2342 -92
rect 2371 -96 2375 -92
rect 359 -290 363 -286
rect 392 -290 396 -286
rect 1102 -293 1106 -289
rect 1135 -293 1139 -289
rect 49 -338 53 -334
rect 82 -338 86 -334
rect 286 -338 290 -334
rect 319 -338 323 -334
rect 1861 -293 1865 -289
rect 1894 -293 1898 -289
rect 792 -341 796 -337
rect 825 -341 829 -337
rect 1029 -341 1033 -337
rect 1062 -341 1066 -337
rect -24 -386 -20 -382
rect 9 -386 13 -382
rect 460 -358 464 -354
rect 493 -358 497 -354
rect 2597 -293 2601 -289
rect 2630 -293 2634 -289
rect 1551 -341 1555 -337
rect 1584 -341 1588 -337
rect 1788 -341 1792 -337
rect 1821 -341 1825 -337
rect 719 -389 723 -385
rect 752 -389 756 -385
rect 374 -399 378 -395
rect 150 -406 154 -402
rect 407 -399 411 -395
rect 183 -406 187 -402
rect 1203 -361 1207 -357
rect 1236 -361 1240 -357
rect 2287 -341 2291 -337
rect 2320 -341 2324 -337
rect 2524 -341 2528 -337
rect 2557 -341 2561 -337
rect 1478 -389 1482 -385
rect 1511 -389 1515 -385
rect 1117 -402 1121 -398
rect 64 -447 68 -443
rect 97 -447 101 -443
rect 893 -409 897 -405
rect 1150 -402 1154 -398
rect 926 -409 930 -405
rect 1962 -361 1966 -357
rect 1995 -361 1999 -357
rect 2214 -389 2218 -385
rect 2247 -389 2251 -385
rect 1876 -402 1880 -398
rect 1652 -409 1656 -405
rect 1909 -402 1913 -398
rect 1685 -409 1689 -405
rect 2698 -361 2702 -357
rect 2731 -361 2735 -357
rect 2612 -402 2616 -398
rect 2388 -409 2392 -405
rect 2645 -402 2649 -398
rect 2421 -409 2425 -405
rect 807 -450 811 -446
rect 840 -450 844 -446
rect 1566 -450 1570 -446
rect 1599 -450 1603 -446
rect 2302 -450 2306 -446
rect 2335 -450 2339 -446
rect 346 -505 350 -501
rect 379 -505 383 -501
rect 412 -505 416 -501
rect 422 -505 426 -501
rect 505 -508 509 -504
rect 515 -508 519 -504
rect 538 -508 542 -504
rect 573 -508 577 -504
rect 583 -508 587 -504
rect 1089 -508 1093 -504
rect 1122 -508 1126 -504
rect 1155 -508 1159 -504
rect 1165 -508 1169 -504
rect 1248 -511 1252 -507
rect 1258 -511 1262 -507
rect 1281 -511 1285 -507
rect 1316 -511 1320 -507
rect 1326 -511 1330 -507
rect 1848 -508 1852 -504
rect 1881 -508 1885 -504
rect 1914 -508 1918 -504
rect 1924 -508 1928 -504
rect 2007 -511 2011 -507
rect 2017 -511 2021 -507
rect 2040 -511 2044 -507
rect 2075 -511 2079 -507
rect 2085 -511 2089 -507
rect 2584 -508 2588 -504
rect 2617 -508 2621 -504
rect 2650 -508 2654 -504
rect 2660 -508 2664 -504
rect 2743 -511 2747 -507
rect 2753 -511 2757 -507
rect 2776 -511 2780 -507
rect 2811 -511 2815 -507
rect 2821 -511 2825 -507
rect 35 -556 39 -552
rect 68 -556 72 -552
rect 101 -556 105 -552
rect 111 -556 115 -552
rect 778 -559 782 -555
rect 811 -559 815 -555
rect 844 -559 848 -555
rect 854 -559 858 -555
rect 1537 -559 1541 -555
rect 1570 -559 1574 -555
rect 1603 -559 1607 -555
rect 1613 -559 1617 -555
rect 2273 -559 2277 -555
rect 2306 -559 2310 -555
rect 2339 -559 2343 -555
rect 2349 -559 2353 -555
<< pdcontact >>
rect 78 58 82 62
rect 88 58 92 62
rect 111 58 115 62
rect 676 58 680 62
rect 686 58 690 62
rect 709 58 713 62
rect 1555 58 1559 62
rect 1565 58 1569 62
rect 1588 58 1592 62
rect 2323 58 2327 62
rect 2333 58 2337 62
rect 2356 58 2360 62
rect 5 10 9 14
rect 15 10 19 14
rect 38 10 42 14
rect 603 10 607 14
rect 613 10 617 14
rect 636 10 640 14
rect 179 -10 183 -6
rect 189 -10 193 -6
rect 212 -10 216 -6
rect 93 -51 97 -47
rect 103 -51 107 -47
rect 126 -51 130 -47
rect 1482 10 1486 14
rect 1492 10 1496 14
rect 1515 10 1519 14
rect 777 -10 781 -6
rect 787 -10 791 -6
rect 810 -10 814 -6
rect 691 -51 695 -47
rect 701 -51 705 -47
rect 724 -51 728 -47
rect 2250 10 2254 14
rect 2260 10 2264 14
rect 2283 10 2287 14
rect 1656 -10 1660 -6
rect 1666 -10 1670 -6
rect 1689 -10 1693 -6
rect 1570 -51 1574 -47
rect 1580 -51 1584 -47
rect 1603 -51 1607 -47
rect 2424 -10 2428 -6
rect 2434 -10 2438 -6
rect 2457 -10 2461 -6
rect 2338 -51 2342 -47
rect 2348 -51 2352 -47
rect 2371 -51 2375 -47
rect 359 -245 363 -241
rect 369 -245 373 -241
rect 392 -245 396 -241
rect 1102 -248 1106 -244
rect 1112 -248 1116 -244
rect 1135 -248 1139 -244
rect 1861 -248 1865 -244
rect 1871 -248 1875 -244
rect 1894 -248 1898 -244
rect 2597 -248 2601 -244
rect 2607 -248 2611 -244
rect 2630 -248 2634 -244
rect 49 -293 53 -289
rect 59 -293 63 -289
rect 82 -293 86 -289
rect 286 -293 290 -289
rect 296 -293 300 -289
rect 319 -293 323 -289
rect 792 -296 796 -292
rect 802 -296 806 -292
rect 825 -296 829 -292
rect 1029 -296 1033 -292
rect 1039 -296 1043 -292
rect 1062 -296 1066 -292
rect 460 -313 464 -309
rect 470 -313 474 -309
rect 493 -313 497 -309
rect -24 -341 -20 -337
rect -14 -341 -10 -337
rect 9 -341 13 -337
rect 374 -354 378 -350
rect 150 -361 154 -357
rect 160 -361 164 -357
rect 384 -354 388 -350
rect 407 -354 411 -350
rect 1551 -296 1555 -292
rect 1561 -296 1565 -292
rect 1584 -296 1588 -292
rect 1788 -296 1792 -292
rect 1798 -296 1802 -292
rect 1821 -296 1825 -292
rect 1203 -316 1207 -312
rect 1213 -316 1217 -312
rect 1236 -316 1240 -312
rect 719 -344 723 -340
rect 729 -344 733 -340
rect 752 -344 756 -340
rect 183 -361 187 -357
rect 64 -402 68 -398
rect 74 -402 78 -398
rect 97 -402 101 -398
rect 1117 -357 1121 -353
rect 893 -364 897 -360
rect 903 -364 907 -360
rect 1127 -357 1131 -353
rect 1150 -357 1154 -353
rect 2287 -296 2291 -292
rect 2297 -296 2301 -292
rect 2320 -296 2324 -292
rect 2524 -296 2528 -292
rect 2534 -296 2538 -292
rect 2557 -296 2561 -292
rect 1962 -316 1966 -312
rect 1972 -316 1976 -312
rect 1995 -316 1999 -312
rect 1478 -344 1482 -340
rect 1488 -344 1492 -340
rect 1511 -344 1515 -340
rect 926 -364 930 -360
rect 807 -405 811 -401
rect 817 -405 821 -401
rect 840 -405 844 -401
rect 1876 -357 1880 -353
rect 1652 -364 1656 -360
rect 1662 -364 1666 -360
rect 1886 -357 1890 -353
rect 1909 -357 1913 -353
rect 2698 -316 2702 -312
rect 2708 -316 2712 -312
rect 2731 -316 2735 -312
rect 2214 -344 2218 -340
rect 2224 -344 2228 -340
rect 2247 -344 2251 -340
rect 1685 -364 1689 -360
rect 1566 -405 1570 -401
rect 1576 -405 1580 -401
rect 1599 -405 1603 -401
rect 2612 -357 2616 -353
rect 2388 -364 2392 -360
rect 2398 -364 2402 -360
rect 2622 -357 2626 -353
rect 2645 -357 2649 -353
rect 2421 -364 2425 -360
rect 2302 -405 2306 -401
rect 2312 -405 2316 -401
rect 2335 -405 2339 -401
rect 346 -460 350 -456
rect 356 -460 360 -456
rect 379 -460 383 -456
rect 412 -460 416 -456
rect 422 -460 426 -456
rect 505 -460 509 -456
rect 540 -460 544 -456
rect 573 -460 577 -456
rect 583 -460 587 -456
rect 35 -511 39 -507
rect 45 -511 49 -507
rect 68 -511 72 -507
rect 101 -511 105 -507
rect 1089 -463 1093 -459
rect 1099 -463 1103 -459
rect 1122 -463 1126 -459
rect 1155 -463 1159 -459
rect 1165 -463 1169 -459
rect 1248 -463 1252 -459
rect 1283 -463 1287 -459
rect 1316 -463 1320 -459
rect 1326 -463 1330 -459
rect 1848 -463 1852 -459
rect 1858 -463 1862 -459
rect 1881 -463 1885 -459
rect 1914 -463 1918 -459
rect 1924 -463 1928 -459
rect 2007 -463 2011 -459
rect 2042 -463 2046 -459
rect 2075 -463 2079 -459
rect 2085 -463 2089 -459
rect 2584 -463 2588 -459
rect 2594 -463 2598 -459
rect 2617 -463 2621 -459
rect 2650 -463 2654 -459
rect 2660 -463 2664 -459
rect 2743 -463 2747 -459
rect 2778 -463 2782 -459
rect 2811 -463 2815 -459
rect 2821 -463 2825 -459
rect 111 -511 115 -507
rect 778 -514 782 -510
rect 788 -514 792 -510
rect 811 -514 815 -510
rect 844 -514 848 -510
rect 854 -514 858 -510
rect 1537 -514 1541 -510
rect 1547 -514 1551 -510
rect 1570 -514 1574 -510
rect 1603 -514 1607 -510
rect 1613 -514 1617 -510
rect 2273 -514 2277 -510
rect 2283 -514 2287 -510
rect 2306 -514 2310 -510
rect 2339 -514 2343 -510
rect 2349 -514 2353 -510
<< polysilicon >>
rect 83 64 87 67
rect 104 64 108 67
rect 681 64 685 67
rect 702 64 706 67
rect 1560 64 1564 67
rect 1581 64 1585 67
rect 2328 64 2332 67
rect 2349 64 2353 67
rect 83 19 87 56
rect 104 19 108 56
rect 681 19 685 56
rect 702 19 706 56
rect 1560 19 1564 56
rect 1581 19 1585 56
rect 2328 19 2332 56
rect 2349 19 2353 56
rect 10 16 14 19
rect 31 16 35 19
rect 608 16 612 19
rect 629 16 633 19
rect 83 8 87 11
rect 10 -29 14 8
rect 31 -29 35 8
rect 104 4 108 11
rect 1487 16 1491 19
rect 1508 16 1512 19
rect 681 8 685 11
rect 184 -4 188 -1
rect 205 -4 209 -1
rect 10 -40 14 -37
rect 31 -45 35 -37
rect 98 -45 102 -42
rect 119 -45 123 -42
rect 184 -49 188 -12
rect 205 -49 209 -12
rect 608 -29 612 8
rect 629 -29 633 8
rect 702 4 706 11
rect 2255 16 2259 19
rect 2276 16 2280 19
rect 1560 8 1564 11
rect 782 -4 786 -1
rect 803 -4 807 -1
rect 608 -40 612 -37
rect 629 -45 633 -37
rect 696 -45 700 -42
rect 717 -45 721 -42
rect 98 -90 102 -53
rect 119 -90 123 -53
rect 782 -49 786 -12
rect 803 -49 807 -12
rect 1487 -29 1491 8
rect 1508 -29 1512 8
rect 1581 4 1585 11
rect 2328 8 2332 11
rect 1661 -4 1665 -1
rect 1682 -4 1686 -1
rect 1487 -40 1491 -37
rect 1508 -45 1512 -37
rect 1575 -45 1579 -42
rect 1596 -45 1600 -42
rect 184 -60 188 -57
rect 205 -65 209 -57
rect 696 -90 700 -53
rect 717 -90 721 -53
rect 1661 -49 1665 -12
rect 1682 -49 1686 -12
rect 2255 -29 2259 8
rect 2276 -29 2280 8
rect 2349 4 2353 11
rect 2429 -4 2433 -1
rect 2450 -4 2454 -1
rect 2255 -40 2259 -37
rect 2276 -45 2280 -37
rect 2343 -45 2347 -42
rect 2364 -45 2368 -42
rect 782 -60 786 -57
rect 803 -65 807 -57
rect 1575 -90 1579 -53
rect 1596 -90 1600 -53
rect 2429 -49 2433 -12
rect 2450 -49 2454 -12
rect 1661 -60 1665 -57
rect 1682 -65 1686 -57
rect 2343 -90 2347 -53
rect 2364 -90 2368 -53
rect 2429 -60 2433 -57
rect 2450 -65 2454 -57
rect 98 -101 102 -98
rect 119 -106 123 -98
rect 696 -101 700 -98
rect 717 -106 721 -98
rect 1575 -101 1579 -98
rect 1596 -106 1600 -98
rect 2343 -101 2347 -98
rect 2364 -106 2368 -98
rect 364 -239 368 -236
rect 385 -239 389 -236
rect 1107 -242 1111 -239
rect 1128 -242 1132 -239
rect 1866 -242 1870 -239
rect 1887 -242 1891 -239
rect 2602 -242 2606 -239
rect 2623 -242 2627 -239
rect 364 -284 368 -247
rect 385 -284 389 -247
rect 54 -287 58 -284
rect 75 -287 79 -284
rect 291 -287 295 -284
rect 312 -287 316 -284
rect 1107 -287 1111 -250
rect 1128 -287 1132 -250
rect 1866 -287 1870 -250
rect 1887 -287 1891 -250
rect 2602 -287 2606 -250
rect 2623 -287 2627 -250
rect 797 -290 801 -287
rect 818 -290 822 -287
rect 1034 -290 1038 -287
rect 1055 -290 1059 -287
rect 364 -295 368 -292
rect 54 -332 58 -295
rect 75 -332 79 -295
rect 291 -332 295 -295
rect 312 -332 316 -295
rect 385 -299 389 -292
rect 1556 -290 1560 -287
rect 1577 -290 1581 -287
rect 1793 -290 1797 -287
rect 1814 -290 1818 -287
rect 1107 -298 1111 -295
rect 465 -307 469 -304
rect 486 -307 490 -304
rect -19 -335 -15 -332
rect 2 -335 6 -332
rect 54 -343 58 -340
rect -19 -380 -15 -343
rect 2 -380 6 -343
rect 75 -347 79 -340
rect 291 -343 295 -340
rect 312 -348 316 -340
rect 379 -348 383 -345
rect 400 -348 404 -345
rect 155 -355 159 -352
rect 176 -355 180 -352
rect 465 -352 469 -315
rect 486 -352 490 -315
rect 797 -335 801 -298
rect 818 -335 822 -298
rect 1034 -335 1038 -298
rect 1055 -335 1059 -298
rect 1128 -302 1132 -295
rect 2292 -290 2296 -287
rect 2313 -290 2317 -287
rect 2529 -290 2533 -287
rect 2550 -290 2554 -287
rect 1866 -298 1870 -295
rect 1208 -310 1212 -307
rect 1229 -310 1233 -307
rect 724 -338 728 -335
rect 745 -338 749 -335
rect 797 -346 801 -343
rect -19 -391 -15 -388
rect 2 -396 6 -388
rect 69 -396 73 -393
rect 90 -396 94 -393
rect 155 -400 159 -363
rect 176 -400 180 -363
rect 379 -393 383 -356
rect 400 -393 404 -356
rect 465 -363 469 -360
rect 486 -368 490 -360
rect 724 -383 728 -346
rect 745 -383 749 -346
rect 818 -350 822 -343
rect 1034 -346 1038 -343
rect 1055 -351 1059 -343
rect 1122 -351 1126 -348
rect 1143 -351 1147 -348
rect 898 -358 902 -355
rect 919 -358 923 -355
rect 1208 -355 1212 -318
rect 1229 -355 1233 -318
rect 1556 -335 1560 -298
rect 1577 -335 1581 -298
rect 1793 -335 1797 -298
rect 1814 -335 1818 -298
rect 1887 -302 1891 -295
rect 2602 -298 2606 -295
rect 1967 -310 1971 -307
rect 1988 -310 1992 -307
rect 1483 -338 1487 -335
rect 1504 -338 1508 -335
rect 1556 -346 1560 -343
rect 69 -441 73 -404
rect 90 -441 94 -404
rect 724 -394 728 -391
rect 745 -399 749 -391
rect 812 -399 816 -396
rect 833 -399 837 -396
rect 379 -404 383 -401
rect 155 -411 159 -408
rect 176 -416 180 -408
rect 400 -409 404 -401
rect 898 -403 902 -366
rect 919 -403 923 -366
rect 1122 -396 1126 -359
rect 1143 -396 1147 -359
rect 1208 -366 1212 -363
rect 1229 -371 1233 -363
rect 1483 -383 1487 -346
rect 1504 -383 1508 -346
rect 1577 -350 1581 -343
rect 1793 -346 1797 -343
rect 1814 -351 1818 -343
rect 1881 -351 1885 -348
rect 1902 -351 1906 -348
rect 1657 -358 1661 -355
rect 1678 -358 1682 -355
rect 1967 -355 1971 -318
rect 1988 -355 1992 -318
rect 2292 -335 2296 -298
rect 2313 -335 2317 -298
rect 2529 -335 2533 -298
rect 2550 -335 2554 -298
rect 2623 -302 2627 -295
rect 2703 -310 2707 -307
rect 2724 -310 2728 -307
rect 2219 -338 2223 -335
rect 2240 -338 2244 -335
rect 2292 -346 2296 -343
rect 1483 -394 1487 -391
rect 812 -444 816 -407
rect 833 -444 837 -407
rect 1504 -399 1508 -391
rect 1571 -399 1575 -396
rect 1592 -399 1596 -396
rect 1122 -407 1126 -404
rect 898 -414 902 -411
rect 919 -419 923 -411
rect 1143 -412 1147 -404
rect 1657 -403 1661 -366
rect 1678 -403 1682 -366
rect 1881 -396 1885 -359
rect 1902 -396 1906 -359
rect 1967 -366 1971 -363
rect 1988 -371 1992 -363
rect 2219 -383 2223 -346
rect 2240 -383 2244 -346
rect 2313 -350 2317 -343
rect 2529 -346 2533 -343
rect 2550 -351 2554 -343
rect 2617 -351 2621 -348
rect 2638 -351 2642 -348
rect 2393 -358 2397 -355
rect 2414 -358 2418 -355
rect 2703 -355 2707 -318
rect 2724 -355 2728 -318
rect 2219 -394 2223 -391
rect 1571 -444 1575 -407
rect 1592 -444 1596 -407
rect 2240 -399 2244 -391
rect 2307 -399 2311 -396
rect 2328 -399 2332 -396
rect 1881 -407 1885 -404
rect 1657 -414 1661 -411
rect 1678 -419 1682 -411
rect 1902 -412 1906 -404
rect 2393 -403 2397 -366
rect 2414 -403 2418 -366
rect 2617 -396 2621 -359
rect 2638 -396 2642 -359
rect 2703 -366 2707 -363
rect 2724 -371 2728 -363
rect 2307 -444 2311 -407
rect 2328 -444 2332 -407
rect 2617 -407 2621 -404
rect 2393 -414 2397 -411
rect 2414 -419 2418 -411
rect 2638 -412 2642 -404
rect 69 -452 73 -449
rect 90 -457 94 -449
rect 351 -454 355 -451
rect 372 -454 376 -451
rect 417 -454 421 -451
rect 510 -454 514 -451
rect 531 -454 535 -451
rect 578 -454 582 -451
rect 812 -455 816 -452
rect 833 -460 837 -452
rect 1094 -457 1098 -454
rect 1115 -457 1119 -454
rect 1160 -457 1164 -454
rect 1253 -457 1257 -454
rect 1274 -457 1278 -454
rect 1321 -457 1325 -454
rect 1571 -455 1575 -452
rect 351 -499 355 -462
rect 372 -499 376 -462
rect 417 -499 421 -462
rect 40 -505 44 -502
rect 61 -505 65 -502
rect 106 -505 110 -502
rect 510 -502 514 -462
rect 531 -502 535 -462
rect 578 -502 582 -462
rect 1592 -460 1596 -452
rect 1853 -457 1857 -454
rect 1874 -457 1878 -454
rect 1919 -457 1923 -454
rect 2012 -457 2016 -454
rect 2033 -457 2037 -454
rect 2080 -457 2084 -454
rect 2307 -455 2311 -452
rect 2328 -460 2332 -452
rect 2589 -457 2593 -454
rect 2610 -457 2614 -454
rect 2655 -457 2659 -454
rect 2748 -457 2752 -454
rect 2769 -457 2773 -454
rect 2816 -457 2820 -454
rect 1094 -502 1098 -465
rect 1115 -502 1119 -465
rect 1160 -502 1164 -465
rect 351 -510 355 -507
rect 372 -510 376 -507
rect 417 -510 421 -507
rect 783 -508 787 -505
rect 804 -508 808 -505
rect 849 -508 853 -505
rect 510 -513 514 -510
rect 531 -513 535 -510
rect 578 -513 582 -510
rect 40 -550 44 -513
rect 61 -550 65 -513
rect 106 -550 110 -513
rect 1253 -505 1257 -465
rect 1274 -505 1278 -465
rect 1321 -505 1325 -465
rect 1853 -502 1857 -465
rect 1874 -502 1878 -465
rect 1919 -502 1923 -465
rect 1094 -513 1098 -510
rect 1115 -513 1119 -510
rect 1160 -513 1164 -510
rect 1542 -508 1546 -505
rect 1563 -508 1567 -505
rect 1608 -508 1612 -505
rect 1253 -516 1257 -513
rect 1274 -516 1278 -513
rect 1321 -516 1325 -513
rect 2012 -505 2016 -465
rect 2033 -505 2037 -465
rect 2080 -505 2084 -465
rect 2589 -502 2593 -465
rect 2610 -502 2614 -465
rect 2655 -502 2659 -465
rect 1853 -513 1857 -510
rect 1874 -513 1878 -510
rect 1919 -513 1923 -510
rect 2278 -508 2282 -505
rect 2299 -508 2303 -505
rect 2344 -508 2348 -505
rect 2012 -516 2016 -513
rect 2033 -516 2037 -513
rect 2080 -516 2084 -513
rect 2748 -505 2752 -465
rect 2769 -505 2773 -465
rect 2816 -505 2820 -465
rect 2589 -513 2593 -510
rect 2610 -513 2614 -510
rect 2655 -513 2659 -510
rect 2748 -516 2752 -513
rect 2769 -516 2773 -513
rect 2816 -516 2820 -513
rect 783 -553 787 -516
rect 804 -553 808 -516
rect 849 -553 853 -516
rect 1542 -553 1546 -516
rect 1563 -553 1567 -516
rect 1608 -553 1612 -516
rect 2278 -553 2282 -516
rect 2299 -553 2303 -516
rect 2344 -553 2348 -516
rect 40 -561 44 -558
rect 61 -561 65 -558
rect 106 -561 110 -558
rect 783 -564 787 -561
rect 804 -564 808 -561
rect 849 -564 853 -561
rect 1542 -564 1546 -561
rect 1563 -564 1567 -561
rect 1608 -564 1612 -561
rect 2278 -564 2282 -561
rect 2299 -564 2303 -561
rect 2344 -564 2348 -561
<< polycontact >>
rect 79 37 83 41
rect 677 37 681 41
rect 1556 37 1560 41
rect 2324 37 2328 41
rect 6 -11 10 -7
rect 100 3 104 7
rect 604 -11 608 -7
rect 180 -31 184 -27
rect 27 -45 31 -41
rect 698 3 702 7
rect 1483 -11 1487 -7
rect 778 -31 782 -27
rect 625 -45 629 -41
rect 94 -72 98 -68
rect 1577 3 1581 7
rect 2251 -11 2255 -7
rect 1657 -31 1661 -27
rect 1504 -45 1508 -41
rect 201 -65 205 -61
rect 692 -72 696 -68
rect 2345 3 2349 7
rect 2425 -31 2429 -27
rect 2272 -45 2276 -41
rect 799 -65 803 -61
rect 1571 -72 1575 -68
rect 1678 -65 1682 -61
rect 2339 -72 2343 -68
rect 2446 -65 2450 -61
rect 115 -106 119 -102
rect 713 -106 717 -102
rect 1592 -106 1596 -102
rect 2360 -106 2364 -102
rect 360 -266 364 -262
rect 1103 -269 1107 -265
rect 1862 -269 1866 -265
rect 2598 -269 2602 -265
rect 50 -314 54 -310
rect 287 -314 291 -310
rect 381 -300 385 -296
rect 461 -334 465 -330
rect -23 -362 -19 -358
rect 71 -348 75 -344
rect 308 -348 312 -344
rect 793 -317 797 -313
rect 1030 -317 1034 -313
rect 1124 -303 1128 -299
rect 1552 -317 1556 -313
rect 1204 -337 1208 -333
rect 151 -382 155 -378
rect -2 -396 2 -392
rect 375 -375 379 -371
rect 482 -368 486 -364
rect 720 -365 724 -361
rect 814 -351 818 -347
rect 1051 -351 1055 -347
rect 1789 -317 1793 -313
rect 1883 -303 1887 -299
rect 2288 -317 2292 -313
rect 1963 -337 1967 -333
rect 894 -385 898 -381
rect 65 -423 69 -419
rect 741 -399 745 -395
rect 172 -416 176 -412
rect 396 -409 400 -405
rect 1118 -378 1122 -374
rect 1225 -371 1229 -367
rect 1479 -365 1483 -361
rect 1573 -351 1577 -347
rect 1810 -351 1814 -347
rect 2525 -317 2529 -313
rect 2619 -303 2623 -299
rect 2699 -337 2703 -333
rect 1653 -385 1657 -381
rect 808 -426 812 -422
rect 1500 -399 1504 -395
rect 915 -419 919 -415
rect 1139 -412 1143 -408
rect 1877 -378 1881 -374
rect 1984 -371 1988 -367
rect 2215 -365 2219 -361
rect 2309 -351 2313 -347
rect 2546 -351 2550 -347
rect 2389 -385 2393 -381
rect 1567 -426 1571 -422
rect 2236 -399 2240 -395
rect 1674 -419 1678 -415
rect 1898 -412 1902 -408
rect 2613 -378 2617 -374
rect 2720 -371 2724 -367
rect 2303 -426 2307 -422
rect 2410 -419 2414 -415
rect 2634 -412 2638 -408
rect 86 -457 90 -453
rect 829 -460 833 -456
rect 347 -481 351 -477
rect 368 -493 372 -489
rect 413 -485 417 -481
rect 506 -482 510 -478
rect 527 -490 531 -486
rect 574 -498 578 -494
rect 1588 -460 1592 -456
rect 2324 -460 2328 -456
rect 1090 -484 1094 -480
rect 1111 -496 1115 -492
rect 1156 -488 1160 -484
rect 1249 -485 1253 -481
rect 36 -532 40 -528
rect 57 -544 61 -540
rect 102 -536 106 -532
rect 1270 -493 1274 -489
rect 1317 -501 1321 -497
rect 1849 -484 1853 -480
rect 1870 -496 1874 -492
rect 1915 -488 1919 -484
rect 2008 -485 2012 -481
rect 2029 -493 2033 -489
rect 2076 -501 2080 -497
rect 2585 -484 2589 -480
rect 2606 -496 2610 -492
rect 2651 -488 2655 -484
rect 2744 -485 2748 -481
rect 2765 -493 2769 -489
rect 2812 -501 2816 -497
rect 779 -535 783 -531
rect 800 -547 804 -543
rect 845 -539 849 -535
rect 1538 -535 1542 -531
rect 1559 -547 1563 -543
rect 1604 -539 1608 -535
rect 2274 -535 2278 -531
rect 2295 -547 2299 -543
rect 2340 -539 2344 -535
<< metal1 >>
rect -76 88 55 92
rect -76 -62 -72 88
rect 51 84 55 88
rect 629 89 644 93
rect 629 84 633 89
rect 47 80 633 84
rect 640 85 644 89
rect 1508 89 1523 93
rect 1508 84 1512 89
rect 645 80 1512 84
rect 1519 85 1523 89
rect 2276 88 2291 92
rect 2276 84 2280 88
rect 1524 80 2280 84
rect 2287 85 2291 88
rect 2292 80 2461 84
rect -14 64 59 68
rect -14 -7 -10 64
rect 55 41 59 64
rect 78 62 82 80
rect 111 62 115 80
rect 55 37 79 41
rect 88 37 92 58
rect 88 33 156 37
rect 5 29 42 33
rect 5 14 9 29
rect 38 14 42 29
rect 111 17 115 33
rect -18 -11 6 -7
rect 15 -11 19 10
rect 96 -11 100 7
rect 15 -15 100 -11
rect 38 -31 42 -15
rect 23 -97 27 -41
rect 68 -68 72 -15
rect 86 -29 134 -25
rect 152 -27 156 33
rect 179 -6 183 80
rect 212 -6 216 80
rect 584 64 657 68
rect 93 -47 97 -29
rect 126 -47 130 -29
rect 152 -31 180 -27
rect 189 -31 193 -10
rect 584 -7 588 64
rect 653 41 657 64
rect 676 62 680 80
rect 709 62 713 80
rect 653 37 677 41
rect 686 37 690 58
rect 686 33 754 37
rect 603 29 640 33
rect 603 14 607 29
rect 636 14 640 29
rect 709 17 713 33
rect 580 -11 604 -7
rect 613 -11 617 10
rect 694 -11 698 7
rect 613 -15 698 -11
rect 636 -31 640 -15
rect 189 -35 237 -31
rect 212 -51 216 -35
rect 68 -72 94 -68
rect 103 -72 107 -51
rect 197 -72 201 -61
rect 621 -68 625 -41
rect 103 -76 201 -72
rect 573 -72 625 -68
rect 666 -68 670 -15
rect 684 -29 732 -25
rect 750 -27 754 33
rect 777 -6 781 80
rect 810 79 1512 80
rect 810 -6 814 79
rect 1463 64 1536 68
rect 691 -47 695 -29
rect 724 -47 728 -29
rect 750 -31 778 -27
rect 787 -31 791 -10
rect 1463 -7 1467 64
rect 1532 41 1536 64
rect 1555 62 1559 80
rect 1588 62 1592 80
rect 1532 37 1556 41
rect 1565 37 1569 58
rect 1565 33 1633 37
rect 1482 29 1519 33
rect 1482 14 1486 29
rect 1515 14 1519 29
rect 1588 17 1592 33
rect 1459 -11 1483 -7
rect 1492 -11 1496 10
rect 1573 -11 1577 7
rect 1492 -15 1577 -11
rect 1515 -31 1519 -15
rect 787 -35 980 -31
rect 810 -51 814 -35
rect 666 -72 692 -68
rect 701 -72 705 -51
rect 795 -72 799 -61
rect 1500 -68 1504 -41
rect 126 -92 130 -76
rect -4 -101 27 -97
rect 23 -121 27 -101
rect 111 -121 115 -102
rect 23 -125 115 -121
rect 573 -129 577 -72
rect 701 -76 799 -72
rect 1453 -76 1504 -68
rect 1545 -68 1549 -15
rect 1563 -29 1611 -25
rect 1629 -27 1633 33
rect 1656 -6 1660 80
rect 1689 -6 1693 80
rect 2218 79 2227 80
rect 2231 64 2304 68
rect 1570 -47 1574 -29
rect 1603 -47 1607 -29
rect 1629 -31 1657 -27
rect 1666 -31 1670 -10
rect 2231 -7 2235 64
rect 2300 41 2304 64
rect 2323 62 2327 80
rect 2356 62 2360 80
rect 2300 37 2324 41
rect 2333 37 2337 58
rect 2333 33 2401 37
rect 2250 29 2287 33
rect 2250 14 2254 29
rect 2283 14 2287 29
rect 2356 17 2360 33
rect 2227 -11 2251 -7
rect 2260 -11 2264 10
rect 2341 -11 2345 7
rect 2260 -15 2345 -11
rect 2283 -31 2287 -15
rect 1666 -35 1750 -31
rect 1689 -51 1693 -35
rect 1545 -72 1571 -68
rect 1580 -72 1584 -51
rect 1674 -72 1678 -61
rect 2268 -68 2272 -41
rect 1580 -76 1678 -72
rect 2214 -76 2272 -68
rect 2313 -68 2317 -15
rect 2331 -29 2379 -25
rect 2397 -27 2401 33
rect 2424 -6 2428 80
rect 2457 -6 2461 80
rect 2338 -47 2342 -29
rect 2371 -47 2375 -29
rect 2397 -31 2425 -27
rect 2434 -31 2438 -10
rect 2434 -35 2484 -31
rect 2457 -51 2461 -35
rect 2313 -72 2339 -68
rect 2348 -72 2352 -51
rect 2442 -72 2446 -61
rect 2348 -76 2446 -72
rect 724 -92 728 -76
rect 709 -129 713 -102
rect -4 -133 713 -129
rect 1453 -148 1457 -76
rect 1500 -121 1504 -76
rect 1603 -92 1607 -76
rect 1588 -121 1592 -102
rect 1500 -125 1592 -121
rect -4 -152 1457 -148
rect 2214 -165 2218 -76
rect 2268 -121 2272 -76
rect 2371 -92 2375 -76
rect 2356 -121 2360 -102
rect 2268 -125 2360 -121
rect -4 -169 2218 -165
rect 328 -223 528 -219
rect 263 -239 340 -235
rect 18 -271 218 -267
rect -47 -287 30 -283
rect -47 -358 -43 -287
rect 26 -310 30 -287
rect 49 -289 53 -271
rect 82 -289 86 -271
rect 26 -314 50 -310
rect 59 -314 63 -293
rect 59 -318 127 -314
rect -24 -322 13 -318
rect -24 -337 -20 -322
rect 9 -337 13 -322
rect 82 -334 86 -318
rect -141 -362 -23 -358
rect -14 -362 -10 -341
rect 67 -362 71 -344
rect -47 -528 -43 -362
rect -14 -366 71 -362
rect 9 -382 13 -366
rect -6 -419 -2 -392
rect -22 -423 -2 -419
rect 39 -419 43 -366
rect 57 -380 105 -376
rect 123 -378 127 -318
rect 150 -357 154 -271
rect 183 -357 187 -271
rect 64 -398 68 -380
rect 97 -398 101 -380
rect 123 -382 151 -378
rect 160 -384 164 -361
rect 160 -388 203 -384
rect 183 -402 187 -388
rect 39 -423 65 -419
rect 74 -423 78 -402
rect 168 -423 172 -412
rect -6 -472 -2 -423
rect 74 -427 172 -423
rect 97 -443 101 -427
rect 82 -472 86 -453
rect -6 -476 86 -472
rect -2 -478 86 -476
rect 214 -485 218 -271
rect 263 -310 267 -239
rect 336 -262 340 -239
rect 359 -241 363 -223
rect 392 -241 396 -223
rect 336 -266 360 -262
rect 369 -266 373 -245
rect 369 -270 437 -266
rect 286 -274 323 -270
rect 286 -289 290 -274
rect 319 -289 323 -274
rect 392 -286 396 -270
rect 238 -314 287 -310
rect 296 -314 300 -293
rect 377 -314 381 -296
rect 263 -477 267 -314
rect 296 -318 381 -314
rect 319 -334 323 -318
rect 304 -371 308 -344
rect 288 -375 308 -371
rect 349 -371 353 -318
rect 367 -332 415 -328
rect 433 -330 437 -270
rect 460 -309 464 -223
rect 493 -309 497 -223
rect 524 -270 528 -223
rect 1071 -226 1271 -222
rect 1830 -226 2030 -222
rect 2566 -226 2766 -222
rect 1006 -242 1083 -238
rect 524 -274 756 -270
rect 761 -274 961 -270
rect 374 -350 378 -332
rect 407 -350 411 -332
rect 433 -334 461 -330
rect 470 -334 474 -313
rect 470 -338 513 -334
rect 493 -354 497 -338
rect 349 -375 375 -371
rect 384 -375 388 -354
rect 478 -375 482 -364
rect 304 -424 308 -375
rect 384 -379 482 -375
rect 407 -395 411 -379
rect 392 -424 396 -405
rect 304 -428 396 -424
rect 524 -434 528 -274
rect 696 -290 773 -286
rect 696 -361 700 -290
rect 769 -313 773 -290
rect 792 -292 796 -274
rect 825 -292 829 -274
rect 769 -317 793 -313
rect 802 -317 806 -296
rect 802 -321 870 -317
rect 719 -325 756 -321
rect 719 -340 723 -325
rect 752 -340 756 -325
rect 825 -337 829 -321
rect 653 -365 720 -361
rect 729 -365 733 -344
rect 810 -365 814 -347
rect 346 -438 577 -434
rect 346 -456 350 -438
rect 379 -456 383 -438
rect 412 -456 416 -438
rect 505 -456 509 -438
rect 573 -456 577 -438
rect 263 -481 347 -477
rect 356 -481 360 -460
rect 422 -478 426 -460
rect 356 -485 413 -481
rect 422 -482 506 -478
rect 35 -489 218 -485
rect 35 -507 39 -489
rect 68 -507 72 -489
rect 101 -507 105 -489
rect 329 -493 368 -489
rect 379 -501 383 -485
rect 422 -501 426 -482
rect 502 -490 527 -486
rect 540 -494 544 -460
rect 583 -481 587 -460
rect 653 -481 657 -365
rect 583 -485 657 -481
rect 515 -498 574 -494
rect 515 -504 519 -498
rect 583 -504 587 -485
rect -47 -532 36 -528
rect 45 -532 49 -511
rect 45 -536 102 -532
rect 19 -544 57 -540
rect 68 -552 72 -536
rect 111 -537 115 -511
rect 346 -520 350 -505
rect 412 -520 416 -505
rect 505 -520 509 -508
rect 538 -520 542 -508
rect 573 -520 577 -508
rect 339 -524 577 -520
rect 111 -541 438 -537
rect 111 -552 115 -541
rect 35 -568 39 -556
rect 101 -568 105 -556
rect 35 -572 105 -568
rect 573 -571 577 -524
rect 696 -531 700 -365
rect 729 -369 814 -365
rect 752 -385 756 -369
rect 737 -422 741 -395
rect 721 -426 741 -422
rect 782 -422 786 -369
rect 800 -383 848 -379
rect 866 -381 870 -321
rect 893 -360 897 -274
rect 926 -360 930 -274
rect 807 -401 811 -383
rect 840 -401 844 -383
rect 866 -385 894 -381
rect 903 -387 907 -364
rect 903 -391 946 -387
rect 926 -405 930 -391
rect 782 -426 808 -422
rect 817 -426 821 -405
rect 911 -426 915 -415
rect 737 -475 741 -426
rect 817 -430 915 -426
rect 840 -446 844 -430
rect 825 -475 829 -456
rect 737 -479 829 -475
rect 957 -488 961 -274
rect 1006 -313 1010 -242
rect 1079 -265 1083 -242
rect 1102 -244 1106 -226
rect 1135 -244 1139 -226
rect 1079 -269 1103 -265
rect 1112 -269 1116 -248
rect 1112 -273 1180 -269
rect 1029 -277 1066 -273
rect 1029 -292 1033 -277
rect 1062 -292 1066 -277
rect 1135 -289 1139 -273
rect 981 -317 1030 -313
rect 1039 -317 1043 -296
rect 1120 -317 1124 -299
rect 1006 -480 1010 -317
rect 1039 -321 1124 -317
rect 1062 -337 1066 -321
rect 1047 -374 1051 -347
rect 1031 -378 1051 -374
rect 1092 -374 1096 -321
rect 1110 -335 1158 -331
rect 1176 -333 1180 -273
rect 1203 -312 1207 -226
rect 1236 -312 1240 -226
rect 1267 -270 1271 -226
rect 1765 -242 1842 -238
rect 1267 -274 1515 -270
rect 1520 -274 1720 -270
rect 1117 -353 1121 -335
rect 1150 -353 1154 -335
rect 1176 -337 1204 -333
rect 1213 -337 1217 -316
rect 1213 -341 1256 -337
rect 1236 -357 1240 -341
rect 1092 -378 1118 -374
rect 1127 -378 1131 -357
rect 1221 -378 1225 -367
rect 1047 -427 1051 -378
rect 1127 -382 1225 -378
rect 1150 -398 1154 -382
rect 1135 -427 1139 -408
rect 1047 -431 1139 -427
rect 1267 -437 1271 -274
rect 1455 -290 1532 -286
rect 1455 -361 1459 -290
rect 1528 -313 1532 -290
rect 1551 -292 1555 -274
rect 1584 -292 1588 -274
rect 1528 -317 1552 -313
rect 1561 -317 1565 -296
rect 1561 -321 1629 -317
rect 1478 -325 1515 -321
rect 1478 -340 1482 -325
rect 1511 -340 1515 -325
rect 1584 -337 1588 -321
rect 1406 -365 1479 -361
rect 1488 -365 1492 -344
rect 1569 -365 1573 -347
rect 1089 -441 1320 -437
rect 1089 -459 1093 -441
rect 1122 -459 1126 -441
rect 1155 -459 1159 -441
rect 1248 -459 1252 -441
rect 1316 -459 1320 -441
rect 1006 -484 1090 -480
rect 1099 -484 1103 -463
rect 1165 -481 1169 -463
rect 1099 -488 1156 -484
rect 1165 -485 1249 -481
rect 778 -492 961 -488
rect 778 -510 782 -492
rect 811 -510 815 -492
rect 844 -510 848 -492
rect 1072 -496 1111 -492
rect 1122 -504 1126 -488
rect 1165 -504 1169 -485
rect 1245 -493 1270 -489
rect 1283 -497 1287 -463
rect 1326 -484 1330 -463
rect 1406 -484 1410 -365
rect 1326 -488 1410 -484
rect 1258 -501 1317 -497
rect 1258 -507 1262 -501
rect 1326 -507 1330 -488
rect 696 -535 779 -531
rect 788 -535 792 -514
rect 788 -539 845 -535
rect 762 -547 800 -543
rect 811 -555 815 -539
rect 854 -540 858 -514
rect 1089 -523 1093 -508
rect 1155 -523 1159 -508
rect 1248 -523 1252 -511
rect 1281 -523 1285 -511
rect 1316 -523 1320 -511
rect 1082 -527 1320 -523
rect 854 -544 1181 -540
rect 854 -555 858 -544
rect 778 -571 782 -559
rect 844 -571 848 -559
rect 1316 -570 1320 -527
rect 1455 -531 1459 -365
rect 1488 -369 1573 -365
rect 1511 -385 1515 -369
rect 1496 -422 1500 -395
rect 1480 -426 1500 -422
rect 1541 -422 1545 -369
rect 1559 -383 1607 -379
rect 1625 -381 1629 -321
rect 1652 -360 1656 -274
rect 1685 -360 1689 -274
rect 1566 -401 1570 -383
rect 1599 -401 1603 -383
rect 1625 -385 1653 -381
rect 1662 -387 1666 -364
rect 1662 -391 1705 -387
rect 1685 -405 1689 -391
rect 1541 -426 1567 -422
rect 1576 -426 1580 -405
rect 1670 -426 1674 -415
rect 1496 -475 1500 -426
rect 1576 -430 1674 -426
rect 1599 -446 1603 -430
rect 1584 -475 1588 -456
rect 1496 -479 1588 -475
rect 1500 -481 1588 -479
rect 1716 -488 1720 -274
rect 1765 -313 1769 -242
rect 1838 -265 1842 -242
rect 1861 -244 1865 -226
rect 1894 -244 1898 -226
rect 1838 -269 1862 -265
rect 1871 -269 1875 -248
rect 1871 -273 1939 -269
rect 1788 -277 1825 -273
rect 1788 -292 1792 -277
rect 1821 -292 1825 -277
rect 1894 -289 1898 -273
rect 1765 -317 1789 -313
rect 1798 -317 1802 -296
rect 1879 -317 1883 -299
rect 1765 -480 1769 -317
rect 1798 -321 1883 -317
rect 1821 -337 1825 -321
rect 1806 -374 1810 -347
rect 1790 -378 1810 -374
rect 1851 -374 1855 -321
rect 1869 -335 1917 -331
rect 1935 -333 1939 -273
rect 1962 -312 1966 -226
rect 1995 -312 1999 -226
rect 2026 -270 2030 -226
rect 2501 -242 2578 -238
rect 2026 -274 2251 -270
rect 2256 -274 2456 -270
rect 1876 -353 1880 -335
rect 1909 -353 1913 -335
rect 1935 -337 1963 -333
rect 1972 -337 1976 -316
rect 1972 -341 2015 -337
rect 1995 -357 1999 -341
rect 1851 -378 1877 -374
rect 1886 -378 1890 -357
rect 1980 -378 1984 -367
rect 1806 -427 1810 -378
rect 1886 -382 1984 -378
rect 1909 -398 1913 -382
rect 2026 -404 2030 -274
rect 2191 -290 2268 -286
rect 2191 -361 2195 -290
rect 2264 -313 2268 -290
rect 2287 -292 2291 -274
rect 2320 -292 2324 -274
rect 2264 -317 2288 -313
rect 2297 -317 2301 -296
rect 2297 -321 2365 -317
rect 2214 -325 2251 -321
rect 2214 -340 2218 -325
rect 2247 -340 2251 -325
rect 2320 -337 2324 -321
rect 2000 -408 2030 -404
rect 2136 -365 2215 -361
rect 2224 -365 2228 -344
rect 2305 -365 2309 -347
rect 1894 -427 1898 -408
rect 1806 -431 1898 -427
rect 2000 -437 2004 -408
rect 1848 -441 2079 -437
rect 1848 -459 1852 -441
rect 1881 -459 1885 -441
rect 1914 -459 1918 -441
rect 2007 -459 2011 -441
rect 2075 -459 2079 -441
rect 1765 -484 1849 -480
rect 1858 -484 1862 -463
rect 1924 -481 1928 -463
rect 1858 -488 1915 -484
rect 1924 -485 2008 -481
rect 1537 -492 1720 -488
rect 1537 -510 1541 -492
rect 1570 -510 1574 -492
rect 1603 -510 1607 -492
rect 1831 -496 1870 -492
rect 1881 -504 1885 -488
rect 1924 -504 1928 -485
rect 2004 -493 2029 -489
rect 2042 -497 2046 -463
rect 2085 -484 2089 -463
rect 2136 -484 2140 -365
rect 2085 -488 2140 -484
rect 2017 -501 2076 -497
rect 2017 -507 2021 -501
rect 2085 -507 2089 -488
rect 1455 -535 1538 -531
rect 1547 -535 1551 -514
rect 1547 -539 1604 -535
rect 1521 -547 1559 -543
rect 1570 -555 1574 -539
rect 1613 -540 1617 -514
rect 1848 -523 1852 -508
rect 1914 -523 1918 -508
rect 2007 -523 2011 -511
rect 2040 -523 2044 -511
rect 2075 -523 2079 -511
rect 1841 -527 2079 -523
rect 1613 -544 1940 -540
rect 1613 -555 1617 -544
rect 1537 -570 1541 -559
rect 1603 -569 1607 -559
rect 573 -575 848 -571
rect 1316 -574 1602 -570
rect 2075 -570 2079 -527
rect 2191 -531 2195 -365
rect 2224 -369 2309 -365
rect 2247 -385 2251 -369
rect 2232 -422 2236 -395
rect 2216 -426 2236 -422
rect 2277 -422 2281 -369
rect 2295 -383 2343 -379
rect 2361 -381 2365 -321
rect 2388 -360 2392 -274
rect 2421 -360 2425 -274
rect 2302 -401 2306 -383
rect 2335 -401 2339 -383
rect 2361 -385 2389 -381
rect 2398 -387 2402 -364
rect 2398 -391 2441 -387
rect 2421 -405 2425 -391
rect 2277 -426 2303 -422
rect 2312 -426 2316 -405
rect 2406 -426 2410 -415
rect 2232 -475 2236 -426
rect 2312 -430 2410 -426
rect 2335 -446 2339 -430
rect 2320 -475 2324 -456
rect 2232 -479 2324 -475
rect 2236 -481 2324 -479
rect 2452 -488 2456 -274
rect 2501 -313 2505 -242
rect 2574 -265 2578 -242
rect 2597 -244 2601 -226
rect 2630 -244 2634 -226
rect 2574 -269 2598 -265
rect 2607 -269 2611 -248
rect 2607 -273 2675 -269
rect 2524 -277 2561 -273
rect 2524 -292 2528 -277
rect 2557 -292 2561 -277
rect 2630 -289 2634 -273
rect 2501 -317 2525 -313
rect 2534 -317 2538 -296
rect 2615 -317 2619 -299
rect 2501 -480 2505 -317
rect 2534 -321 2619 -317
rect 2557 -337 2561 -321
rect 2542 -374 2546 -347
rect 2526 -378 2546 -374
rect 2587 -374 2591 -321
rect 2605 -335 2653 -331
rect 2671 -333 2675 -273
rect 2698 -312 2702 -226
rect 2731 -312 2735 -226
rect 2612 -353 2616 -335
rect 2645 -353 2649 -335
rect 2671 -337 2699 -333
rect 2708 -337 2712 -316
rect 2708 -341 2751 -337
rect 2731 -357 2735 -341
rect 2587 -378 2613 -374
rect 2622 -378 2626 -357
rect 2716 -378 2720 -367
rect 2542 -427 2546 -378
rect 2622 -382 2720 -378
rect 2645 -398 2649 -382
rect 2762 -404 2766 -226
rect 2736 -408 2766 -404
rect 2630 -427 2634 -408
rect 2542 -431 2634 -427
rect 2736 -437 2740 -408
rect 2584 -441 2815 -437
rect 2584 -459 2588 -441
rect 2617 -459 2621 -441
rect 2650 -459 2654 -441
rect 2743 -459 2747 -441
rect 2811 -459 2815 -441
rect 2501 -484 2585 -480
rect 2594 -484 2598 -463
rect 2660 -481 2664 -463
rect 2594 -488 2651 -484
rect 2660 -485 2744 -481
rect 2273 -492 2456 -488
rect 2273 -510 2277 -492
rect 2306 -510 2310 -492
rect 2339 -510 2343 -492
rect 2567 -496 2606 -492
rect 2617 -504 2621 -488
rect 2660 -504 2664 -485
rect 2740 -493 2765 -489
rect 2778 -497 2782 -463
rect 2821 -484 2825 -463
rect 2821 -488 2833 -484
rect 2753 -501 2812 -497
rect 2753 -507 2757 -501
rect 2821 -507 2825 -488
rect 2191 -535 2274 -531
rect 2283 -535 2287 -514
rect 2283 -539 2340 -535
rect 2257 -547 2295 -543
rect 2306 -555 2310 -539
rect 2349 -540 2353 -514
rect 2584 -523 2588 -508
rect 2650 -523 2654 -508
rect 2743 -523 2747 -511
rect 2776 -523 2780 -511
rect 2811 -523 2815 -511
rect 2577 -527 2815 -523
rect 2349 -544 2676 -540
rect 2349 -555 2353 -544
rect 2273 -570 2277 -559
rect 2339 -568 2343 -559
rect 2075 -573 2338 -570
rect -141 -626 668 -622
rect 1442 -639 1446 -635
rect -141 -643 1446 -639
rect 2166 -656 2170 -646
rect -141 -660 2170 -656
<< m2contact >>
rect 42 80 47 85
rect 640 80 645 85
rect 1519 80 1524 85
rect 2287 80 2292 85
rect -27 -11 -18 -6
rect 37 33 42 38
rect 77 8 82 13
rect 4 -40 9 -35
rect -77 -68 -72 -62
rect 134 -29 139 -24
rect 174 14 179 19
rect 571 -11 580 -6
rect 635 33 640 38
rect 675 8 680 13
rect 602 -40 607 -35
rect 178 -60 183 -55
rect 732 -29 737 -24
rect 772 14 777 19
rect 1450 -11 1459 -6
rect 1514 33 1519 38
rect 1554 8 1559 13
rect 1481 -40 1486 -35
rect 776 -60 781 -55
rect 92 -101 97 -96
rect 1611 -29 1616 -24
rect 1651 14 1656 19
rect 2218 -11 2227 -6
rect 2282 33 2287 38
rect 2322 8 2327 13
rect 2249 -40 2254 -35
rect 1655 -60 1660 -55
rect 2379 -29 2384 -24
rect 2419 14 2424 19
rect 2423 -60 2428 -55
rect 690 -101 695 -96
rect 1569 -101 1574 -96
rect 2337 -101 2342 -96
rect 323 -223 328 -218
rect 13 -271 18 -266
rect 8 -318 13 -313
rect 48 -343 53 -338
rect -25 -391 -20 -386
rect 105 -380 110 -375
rect 145 -337 150 -332
rect 203 -388 208 -383
rect 149 -411 154 -406
rect -22 -428 -17 -423
rect 63 -452 68 -447
rect 318 -270 323 -265
rect 358 -295 363 -290
rect 285 -343 290 -338
rect 415 -332 420 -327
rect 455 -289 460 -284
rect 1066 -226 1071 -221
rect 1825 -226 1830 -221
rect 2561 -226 2566 -221
rect 756 -274 761 -269
rect 513 -338 518 -333
rect 459 -363 464 -358
rect 288 -380 293 -375
rect 373 -404 378 -399
rect 751 -321 756 -316
rect 791 -346 796 -341
rect 324 -494 329 -489
rect 14 -545 19 -540
rect 340 -530 345 -524
rect 438 -541 443 -536
rect 105 -572 110 -567
rect 718 -394 723 -389
rect 848 -383 853 -378
rect 888 -340 893 -335
rect 946 -391 951 -386
rect 892 -414 897 -409
rect 721 -431 726 -426
rect 806 -455 811 -450
rect 1061 -273 1066 -268
rect 1101 -298 1106 -293
rect 1028 -346 1033 -341
rect 1158 -335 1163 -330
rect 1198 -292 1203 -287
rect 1515 -274 1520 -269
rect 1256 -341 1261 -336
rect 1202 -366 1207 -361
rect 1031 -383 1036 -378
rect 1116 -407 1121 -402
rect 1510 -321 1515 -316
rect 1550 -346 1555 -341
rect 1067 -497 1072 -492
rect 757 -548 762 -543
rect 1083 -533 1088 -527
rect 1181 -544 1186 -539
rect 1477 -394 1482 -389
rect 1607 -383 1612 -378
rect 1647 -340 1652 -335
rect 1705 -391 1710 -386
rect 1651 -414 1656 -409
rect 1480 -431 1485 -426
rect 1565 -455 1570 -450
rect 1820 -273 1825 -268
rect 1860 -298 1865 -293
rect 1787 -346 1792 -341
rect 1917 -335 1922 -330
rect 1957 -292 1962 -287
rect 2251 -274 2256 -269
rect 2015 -341 2020 -336
rect 1961 -366 1966 -361
rect 1790 -383 1795 -378
rect 1875 -407 1880 -402
rect 2246 -321 2251 -316
rect 2286 -346 2291 -341
rect 1826 -497 1831 -492
rect 1516 -548 1521 -543
rect 1842 -533 1847 -527
rect 1940 -544 1945 -539
rect 848 -575 853 -570
rect 1602 -574 1607 -569
rect 2213 -394 2218 -389
rect 2343 -383 2348 -378
rect 2383 -340 2388 -335
rect 2441 -391 2446 -386
rect 2387 -414 2392 -409
rect 2216 -431 2221 -426
rect 2301 -455 2306 -450
rect 2556 -273 2561 -268
rect 2596 -298 2601 -293
rect 2523 -346 2528 -341
rect 2653 -335 2658 -330
rect 2693 -292 2698 -287
rect 2751 -341 2756 -336
rect 2697 -366 2702 -361
rect 2526 -383 2531 -378
rect 2611 -407 2616 -402
rect 2562 -497 2567 -492
rect 2252 -548 2257 -543
rect 2578 -533 2583 -527
rect 2676 -544 2681 -539
rect 2338 -573 2343 -568
rect 668 -626 673 -621
rect 1441 -635 1446 -630
rect 2166 -646 2171 -641
<< pdm12contact >>
rect 497 -490 502 -485
rect 1240 -493 1245 -488
rect 1999 -493 2004 -488
rect 2735 -493 2740 -488
<< metal2 >>
rect -27 99 -23 107
rect -131 95 2226 99
rect -131 -432 -127 95
rect -27 -6 -23 95
rect 38 38 42 84
rect 139 14 174 18
rect 5 -49 9 -40
rect 78 -49 82 8
rect 139 -29 143 14
rect 571 -6 575 95
rect 636 38 640 84
rect 737 14 772 18
rect 603 -49 607 -40
rect 676 -49 680 8
rect 737 -29 741 14
rect 1450 -6 1458 95
rect 1515 38 1519 84
rect 1616 14 1651 18
rect 1482 -49 1486 -40
rect 1555 -49 1559 8
rect 1616 -29 1620 14
rect 2218 -6 2226 95
rect 2283 38 2287 84
rect 2384 14 2419 18
rect 2250 -49 2254 -40
rect 2323 -49 2327 8
rect 2384 -29 2388 14
rect -120 -53 82 -49
rect 596 -53 680 -49
rect 1475 -53 1559 -49
rect 2243 -53 2327 -49
rect -120 -400 -116 -53
rect -76 -219 -72 -68
rect 78 -110 82 -53
rect 93 -110 97 -101
rect 179 -110 183 -60
rect 676 -110 680 -53
rect 691 -110 695 -101
rect 777 -110 781 -60
rect 1555 -110 1559 -53
rect 1570 -110 1574 -101
rect 1656 -110 1660 -60
rect 2323 -110 2327 -53
rect 2338 -110 2342 -101
rect 2424 -110 2428 -60
rect 78 -114 2428 -110
rect -76 -223 323 -219
rect 9 -313 13 -223
rect 319 -265 323 -223
rect 752 -226 1066 -222
rect 1511 -226 1825 -222
rect 2247 -226 2561 -222
rect 420 -289 455 -285
rect 110 -337 145 -333
rect -24 -400 -20 -391
rect 49 -400 53 -343
rect 110 -380 114 -337
rect 286 -352 290 -343
rect 359 -352 363 -295
rect 420 -332 424 -289
rect 752 -316 756 -226
rect 1062 -268 1066 -226
rect 1163 -292 1198 -288
rect 518 -338 536 -334
rect 853 -340 888 -336
rect 286 -356 363 -352
rect 289 -384 293 -380
rect 208 -388 293 -384
rect -120 -404 53 -400
rect -21 -432 -17 -428
rect -131 -436 -17 -432
rect -21 -540 -17 -436
rect 49 -461 53 -404
rect 64 -461 68 -452
rect 150 -461 154 -411
rect 49 -465 154 -461
rect -21 -544 14 -540
rect 150 -568 154 -465
rect 289 -489 293 -388
rect 359 -413 363 -356
rect 374 -413 378 -404
rect 460 -413 464 -363
rect 719 -403 723 -394
rect 792 -403 796 -346
rect 853 -383 857 -340
rect 1029 -355 1033 -346
rect 1102 -355 1106 -298
rect 1163 -335 1167 -292
rect 1511 -316 1515 -226
rect 1821 -268 1825 -226
rect 1922 -292 1957 -288
rect 1261 -341 1279 -337
rect 1612 -340 1647 -336
rect 1029 -359 1106 -355
rect 1032 -387 1036 -383
rect 951 -391 1036 -387
rect 712 -407 796 -403
rect 359 -417 464 -413
rect 289 -493 324 -489
rect 460 -526 464 -417
rect 722 -435 726 -431
rect 673 -439 726 -435
rect 345 -530 464 -526
rect 472 -490 497 -486
rect 374 -568 378 -530
rect 472 -536 476 -490
rect 443 -540 476 -536
rect 110 -572 378 -568
rect 673 -626 677 -439
rect 722 -543 726 -439
rect 792 -464 796 -407
rect 807 -464 811 -455
rect 893 -464 897 -414
rect 792 -468 897 -464
rect 722 -547 757 -543
rect 893 -571 897 -468
rect 1032 -492 1036 -391
rect 1102 -416 1106 -359
rect 1117 -416 1121 -407
rect 1203 -416 1207 -366
rect 1478 -403 1482 -394
rect 1551 -403 1555 -346
rect 1612 -383 1616 -340
rect 1788 -355 1792 -346
rect 1861 -355 1865 -298
rect 1922 -335 1926 -292
rect 2247 -316 2251 -226
rect 2557 -268 2561 -226
rect 2658 -292 2693 -288
rect 2020 -341 2036 -337
rect 2348 -340 2383 -336
rect 1788 -359 1865 -355
rect 1791 -387 1795 -383
rect 1710 -391 1795 -387
rect 1478 -407 1555 -403
rect 1102 -420 1207 -416
rect 1032 -496 1067 -492
rect 1203 -529 1207 -420
rect 1481 -435 1485 -431
rect 1442 -439 1485 -435
rect 1088 -533 1207 -529
rect 1215 -493 1240 -489
rect 1117 -571 1121 -533
rect 1215 -539 1219 -493
rect 1186 -543 1219 -539
rect 853 -575 1121 -571
rect 1442 -630 1446 -439
rect 1481 -543 1485 -439
rect 1551 -464 1555 -407
rect 1566 -464 1570 -455
rect 1652 -464 1656 -414
rect 1551 -468 1656 -464
rect 1481 -547 1516 -543
rect 1652 -570 1656 -468
rect 1791 -492 1795 -391
rect 1861 -416 1865 -359
rect 1876 -416 1880 -407
rect 1962 -416 1966 -366
rect 2214 -403 2218 -394
rect 2287 -403 2291 -346
rect 2348 -383 2352 -340
rect 2524 -355 2528 -346
rect 2597 -355 2601 -298
rect 2658 -335 2662 -292
rect 2756 -341 2772 -337
rect 2524 -359 2601 -355
rect 2527 -387 2531 -383
rect 2446 -391 2531 -387
rect 2214 -407 2291 -403
rect 1861 -420 1966 -416
rect 1791 -496 1826 -492
rect 1962 -529 1966 -420
rect 2217 -435 2221 -431
rect 2166 -439 2221 -435
rect 1847 -533 1966 -529
rect 1974 -493 1999 -489
rect 1876 -570 1880 -533
rect 1974 -539 1978 -493
rect 1945 -543 1978 -539
rect 1607 -574 1880 -570
rect 2166 -641 2170 -439
rect 2217 -543 2221 -439
rect 2287 -464 2291 -407
rect 2302 -464 2306 -455
rect 2388 -464 2392 -414
rect 2287 -468 2392 -464
rect 2217 -547 2252 -543
rect 2388 -570 2392 -468
rect 2527 -492 2531 -391
rect 2597 -416 2601 -359
rect 2612 -416 2616 -407
rect 2698 -416 2702 -366
rect 2597 -420 2702 -416
rect 2527 -496 2562 -492
rect 2698 -529 2702 -420
rect 2583 -533 2702 -529
rect 2710 -493 2735 -489
rect 2612 -570 2616 -533
rect 2710 -539 2714 -493
rect 2681 -543 2714 -539
rect 2343 -573 2616 -570
<< m123contact >>
rect 232 -40 237 -35
rect 976 -40 981 -35
rect 1745 -40 1750 -35
rect 2479 -40 2484 -35
rect 233 -314 238 -309
rect 976 -317 981 -312
rect 1760 -317 1765 -312
rect 2496 -317 2501 -312
<< metal3 >>
rect 233 -309 237 -40
rect 976 -312 980 -40
rect 1746 -313 1750 -40
rect 1746 -317 1760 -313
rect 2480 -313 2484 -40
rect 2480 -317 2496 -313
<< labels >>
rlabel metal2 0 -52 4 -51 1 GND
rlabel metal1 51 81 55 82 1 VDD
rlabel metal1 825 -34 828 -33 1 B1new
rlabel metal1 1704 -34 1707 -33 1 B2new
rlabel metal1 -2 -101 1 -99 1 B0
rlabel metal1 -1 -132 4 -130 1 B1
rlabel metal1 -135 -360 -132 -358 3 A0
rlabel metal2 -26 101 -24 102 1 M
rlabel metal1 0 -167 5 -165 1 B3
rlabel metal1 233 -34 236 -33 1 B0new
rlabel metal2 531 -337 534 -336 1 s0
rlabel metal1 -2 -152 3 -150 1 B2
rlabel metal1 -139 -625 -136 -624 3 A1
rlabel metal2 1273 -340 1277 -339 1 s1
rlabel metal1 -139 -643 -134 -641 3 A2
rlabel metal1 -140 -659 -136 -657 2 A3
rlabel metal2 2034 -340 2036 -338 1 s2
rlabel metal1 2470 -34 2473 -33 1 B3new
rlabel metal2 2768 -340 2770 -338 1 s3
rlabel metal1 2826 -487 2828 -486 1 carry
<< end >>
