magic
tech scmos
timestamp 1700496324
<< nwell >>
rect -58 0 -30 24
rect 18 0 78 24
rect 84 0 112 24
rect 184 0 244 24
rect 250 0 278 24
rect -55 -109 -27 -85
rect 18 -109 78 -85
rect 84 -109 112 -85
rect 184 -109 244 -85
rect 250 -109 278 -85
<< ntransistor >>
rect -46 -31 -42 -23
rect 30 -37 34 -29
rect 51 -37 55 -29
rect 96 -37 100 -29
rect 196 -37 200 -29
rect 217 -37 221 -29
rect 262 -37 266 -29
rect -43 -140 -39 -132
rect 30 -146 34 -138
rect 51 -146 55 -138
rect 96 -146 100 -138
rect 196 -146 200 -138
rect 217 -146 221 -138
rect 262 -146 266 -138
<< ptransistor >>
rect -46 8 -42 16
rect 30 8 34 16
rect 51 8 55 16
rect 96 8 100 16
rect 196 8 200 16
rect 217 8 221 16
rect 262 8 266 16
rect -43 -101 -39 -93
rect 30 -101 34 -93
rect 51 -101 55 -93
rect 96 -101 100 -93
rect 196 -101 200 -93
rect 217 -101 221 -93
rect 262 -101 266 -93
<< ndiffusion >>
rect -52 -25 -46 -23
rect -52 -29 -51 -25
rect -47 -29 -46 -25
rect -52 -31 -46 -29
rect -42 -25 -36 -23
rect -42 -29 -41 -25
rect -37 -29 -36 -25
rect -42 -31 -36 -29
rect 24 -31 30 -29
rect 24 -35 25 -31
rect 29 -35 30 -31
rect 24 -37 30 -35
rect 34 -37 51 -29
rect 55 -31 72 -29
rect 55 -35 58 -31
rect 62 -35 72 -31
rect 55 -37 72 -35
rect 90 -31 96 -29
rect 90 -35 91 -31
rect 95 -35 96 -31
rect 90 -37 96 -35
rect 100 -31 106 -29
rect 100 -35 101 -31
rect 105 -35 106 -31
rect 100 -37 106 -35
rect 190 -31 196 -29
rect 190 -35 191 -31
rect 195 -35 196 -31
rect 190 -37 196 -35
rect 200 -37 217 -29
rect 221 -31 238 -29
rect 221 -35 224 -31
rect 228 -35 238 -31
rect 221 -37 238 -35
rect 256 -31 262 -29
rect 256 -35 257 -31
rect 261 -35 262 -31
rect 256 -37 262 -35
rect 266 -31 272 -29
rect 266 -35 267 -31
rect 271 -35 272 -31
rect 266 -37 272 -35
rect -49 -134 -43 -132
rect -49 -138 -48 -134
rect -44 -138 -43 -134
rect -49 -140 -43 -138
rect -39 -134 -33 -132
rect -39 -138 -38 -134
rect -34 -138 -33 -134
rect -39 -140 -33 -138
rect 24 -140 30 -138
rect 24 -144 25 -140
rect 29 -144 30 -140
rect 24 -146 30 -144
rect 34 -146 51 -138
rect 55 -140 72 -138
rect 55 -144 58 -140
rect 62 -144 72 -140
rect 55 -146 72 -144
rect 90 -140 96 -138
rect 90 -144 91 -140
rect 95 -144 96 -140
rect 90 -146 96 -144
rect 100 -140 106 -138
rect 100 -144 101 -140
rect 105 -144 106 -140
rect 100 -146 106 -144
rect 190 -140 196 -138
rect 190 -144 191 -140
rect 195 -144 196 -140
rect 190 -146 196 -144
rect 200 -146 217 -138
rect 221 -140 238 -138
rect 221 -144 224 -140
rect 228 -144 238 -140
rect 221 -146 238 -144
rect 256 -140 262 -138
rect 256 -144 257 -140
rect 261 -144 262 -140
rect 256 -146 262 -144
rect 266 -140 272 -138
rect 266 -144 267 -140
rect 271 -144 272 -140
rect 266 -146 272 -144
<< pdiffusion >>
rect -52 14 -46 16
rect -52 10 -51 14
rect -47 10 -46 14
rect -52 8 -46 10
rect -42 14 -36 16
rect -42 10 -41 14
rect -37 10 -36 14
rect -42 8 -36 10
rect 24 14 30 16
rect 24 10 25 14
rect 29 10 30 14
rect 24 8 30 10
rect 34 14 51 16
rect 34 10 35 14
rect 39 10 51 14
rect 34 8 51 10
rect 55 14 72 16
rect 55 10 58 14
rect 62 10 72 14
rect 55 8 72 10
rect 90 14 96 16
rect 90 10 91 14
rect 95 10 96 14
rect 90 8 96 10
rect 100 14 106 16
rect 100 10 101 14
rect 105 10 106 14
rect 100 8 106 10
rect 190 14 196 16
rect 190 10 191 14
rect 195 10 196 14
rect 190 8 196 10
rect 200 14 217 16
rect 200 10 201 14
rect 205 10 217 14
rect 200 8 217 10
rect 221 14 238 16
rect 221 10 224 14
rect 228 10 238 14
rect 221 8 238 10
rect 256 14 262 16
rect 256 10 257 14
rect 261 10 262 14
rect 256 8 262 10
rect 266 14 272 16
rect 266 10 267 14
rect 271 10 272 14
rect 266 8 272 10
rect -49 -95 -43 -93
rect -49 -99 -48 -95
rect -44 -99 -43 -95
rect -49 -101 -43 -99
rect -39 -95 -33 -93
rect -39 -99 -38 -95
rect -34 -99 -33 -95
rect -39 -101 -33 -99
rect 24 -95 30 -93
rect 24 -99 25 -95
rect 29 -99 30 -95
rect 24 -101 30 -99
rect 34 -95 51 -93
rect 34 -99 35 -95
rect 39 -99 51 -95
rect 34 -101 51 -99
rect 55 -95 72 -93
rect 55 -99 58 -95
rect 62 -99 72 -95
rect 55 -101 72 -99
rect 90 -95 96 -93
rect 90 -99 91 -95
rect 95 -99 96 -95
rect 90 -101 96 -99
rect 100 -95 106 -93
rect 100 -99 101 -95
rect 105 -99 106 -95
rect 100 -101 106 -99
rect 190 -95 196 -93
rect 190 -99 191 -95
rect 195 -99 196 -95
rect 190 -101 196 -99
rect 200 -95 217 -93
rect 200 -99 201 -95
rect 205 -99 217 -95
rect 200 -101 217 -99
rect 221 -95 238 -93
rect 221 -99 224 -95
rect 228 -99 238 -95
rect 221 -101 238 -99
rect 256 -95 262 -93
rect 256 -99 257 -95
rect 261 -99 262 -95
rect 256 -101 262 -99
rect 266 -95 272 -93
rect 266 -99 267 -95
rect 271 -99 272 -95
rect 266 -101 272 -99
<< ndcontact >>
rect -51 -29 -47 -25
rect -41 -29 -37 -25
rect 25 -35 29 -31
rect 58 -35 62 -31
rect 91 -35 95 -31
rect 101 -35 105 -31
rect 191 -35 195 -31
rect 224 -35 228 -31
rect 257 -35 261 -31
rect 267 -35 271 -31
rect -48 -138 -44 -134
rect -38 -138 -34 -134
rect 25 -144 29 -140
rect 58 -144 62 -140
rect 91 -144 95 -140
rect 101 -144 105 -140
rect 191 -144 195 -140
rect 224 -144 228 -140
rect 257 -144 261 -140
rect 267 -144 271 -140
<< pdcontact >>
rect -51 10 -47 14
rect -41 10 -37 14
rect 25 10 29 14
rect 35 10 39 14
rect 58 10 62 14
rect 91 10 95 14
rect 101 10 105 14
rect 191 10 195 14
rect 201 10 205 14
rect 224 10 228 14
rect 257 10 261 14
rect 267 10 271 14
rect -48 -99 -44 -95
rect -38 -99 -34 -95
rect 25 -99 29 -95
rect 35 -99 39 -95
rect 58 -99 62 -95
rect 91 -99 95 -95
rect 101 -99 105 -95
rect 191 -99 195 -95
rect 201 -99 205 -95
rect 224 -99 228 -95
rect 257 -99 261 -95
rect 267 -99 271 -95
<< polysilicon >>
rect -46 16 -42 19
rect 30 16 34 19
rect 51 16 55 19
rect 96 16 100 19
rect 196 16 200 19
rect 217 16 221 19
rect 262 16 266 19
rect -46 -23 -42 8
rect 30 -29 34 8
rect 51 -29 55 8
rect 96 -29 100 8
rect 196 -29 200 8
rect 217 -29 221 8
rect 262 -29 266 8
rect -46 -34 -42 -31
rect 30 -40 34 -37
rect 51 -40 55 -37
rect 96 -40 100 -37
rect 196 -40 200 -37
rect 217 -40 221 -37
rect 262 -40 266 -37
rect -43 -93 -39 -90
rect 30 -93 34 -90
rect 51 -93 55 -90
rect 96 -93 100 -90
rect 196 -93 200 -90
rect 217 -93 221 -90
rect 262 -93 266 -90
rect -43 -132 -39 -101
rect 30 -138 34 -101
rect 51 -138 55 -101
rect 96 -138 100 -101
rect 196 -138 200 -101
rect 217 -138 221 -101
rect 262 -138 266 -101
rect -43 -143 -39 -140
rect 30 -149 34 -146
rect 51 -149 55 -146
rect 96 -149 100 -146
rect 196 -149 200 -146
rect 217 -149 221 -146
rect 262 -149 266 -146
<< polycontact >>
rect -50 -11 -46 -7
rect 26 -11 30 -7
rect 47 -23 51 -19
rect 92 -15 96 -11
rect 192 -11 196 -7
rect 213 -23 217 -19
rect 258 -15 262 -11
rect -47 -120 -43 -116
rect 26 -120 30 -116
rect 47 -132 51 -128
rect 92 -124 96 -120
rect 192 -120 196 -116
rect 213 -132 217 -128
rect 258 -124 262 -120
<< metal1 >>
rect -94 57 173 61
rect -94 -45 -90 57
rect -80 49 158 53
rect -80 -7 -76 49
rect -65 32 104 36
rect -51 14 -47 32
rect 25 14 29 32
rect 58 14 62 32
rect 91 14 95 32
rect -80 -11 -50 -7
rect -41 -11 -37 10
rect 22 -11 26 -7
rect 35 -11 39 10
rect -41 -15 -23 -11
rect 35 -15 92 -11
rect -41 -25 -37 -15
rect -51 -45 -47 -29
rect -94 -49 -47 -45
rect -27 -45 -23 -15
rect 6 -23 47 -19
rect 6 -45 10 -23
rect 58 -31 62 -15
rect 101 -16 105 10
rect 101 -20 135 -16
rect 101 -31 105 -20
rect -27 -49 10 -45
rect 25 -45 29 -35
rect 91 -45 95 -35
rect 25 -49 95 -45
rect -78 -154 -74 -49
rect 6 -64 10 -49
rect -48 -77 104 -73
rect -48 -95 -44 -77
rect 25 -95 29 -77
rect 58 -95 62 -77
rect 91 -95 95 -77
rect -62 -120 -47 -116
rect -38 -120 -34 -99
rect 2 -120 26 -116
rect 35 -120 39 -99
rect -38 -124 -20 -120
rect -38 -134 -34 -124
rect 35 -124 92 -120
rect 11 -132 47 -128
rect -48 -154 -44 -138
rect 58 -140 62 -124
rect 101 -125 105 -99
rect 101 -129 120 -125
rect 101 -140 105 -129
rect 25 -154 29 -144
rect 91 -154 95 -144
rect -78 -158 95 -154
rect 116 -181 120 -129
rect 131 -181 135 -20
rect 154 -19 158 49
rect 169 28 173 57
rect 184 32 261 36
rect 191 14 195 32
rect 224 14 228 32
rect 257 14 261 32
rect 188 -11 192 -7
rect 201 -11 205 10
rect 201 -15 258 -11
rect 154 -23 213 -19
rect 154 -128 158 -23
rect 224 -31 228 -15
rect 267 -16 271 10
rect 267 -20 278 -16
rect 267 -31 271 -20
rect 191 -45 195 -35
rect 257 -45 261 -35
rect 184 -49 261 -45
rect 167 -77 261 -73
rect 191 -95 195 -77
rect 224 -95 228 -77
rect 257 -95 261 -77
rect 188 -120 192 -116
rect 201 -120 205 -99
rect 201 -124 258 -120
rect 154 -132 213 -128
rect 224 -140 228 -124
rect 267 -125 271 -99
rect 267 -129 278 -125
rect 267 -140 271 -129
rect 191 -154 195 -144
rect 257 -154 261 -144
rect 188 -158 261 -154
<< m2contact >>
rect 17 -11 22 -6
rect 5 -69 10 -64
rect -67 -120 -62 -115
rect -3 -120 2 -115
rect -20 -125 -15 -120
rect 6 -132 11 -127
rect 183 -11 188 -6
rect 183 -120 188 -115
<< metal2 >>
rect -11 44 163 48
rect -11 -7 -7 44
rect -11 -11 17 -7
rect 159 -7 163 44
rect 159 -11 183 -7
rect -71 -169 -67 -116
rect -11 -121 -7 -11
rect -15 -125 -7 -121
rect -3 -169 1 -120
rect 6 -127 10 -69
rect 160 -120 183 -116
rect 160 -169 164 -120
rect -71 -173 164 -169
<< m123contact >>
rect -70 32 -65 37
rect 104 32 109 37
rect 179 32 184 37
rect 168 23 173 28
rect -53 -77 -48 -72
rect 95 -49 100 -44
rect 179 -49 184 -44
rect 104 -77 109 -72
rect 162 -77 167 -72
rect 95 -158 100 -153
rect 183 -158 188 -153
<< metal3 >>
rect -86 32 -70 36
rect 109 32 179 36
rect -86 -73 -82 32
rect 169 -45 173 23
rect 100 -49 179 -45
rect 169 -61 173 -49
rect 169 -65 177 -61
rect -86 -77 -53 -73
rect 109 -77 162 -73
rect 173 -154 177 -65
rect 100 -158 183 -154
<< labels >>
rlabel metal1 -62 -11 -58 -8 1 S0
rlabel metal1 -54 34 -52 35 4 VDD
rlabel metal1 -54 -48 -52 -47 2 GND
rlabel metal1 -36 -14 -32 -13 1 S0comp
rlabel metal1 181 -22 185 -21 1 S0
rlabel metal2 175 -10 178 -9 1 S1comp
rlabel metal1 12 -23 16 -22 1 S0comp
rlabel metal2 2 -11 5 -9 1 S1comp
rlabel metal1 -59 -120 -55 -118 1 S1
rlabel metal1 -32 -123 -29 -122 1 S1comp
rlabel metal1 12 -132 16 -131 1 S0comp
rlabel metal1 14 -119 18 -117 1 S1
rlabel metal1 181 -131 185 -130 1 S0
rlabel metal2 179 -119 182 -118 1 S1
rlabel metal1 117 -180 119 -179 1 D2
rlabel metal1 132 -180 134 -179 1 D0
rlabel metal1 274 -128 277 -127 7 D3
rlabel metal1 275 -19 278 -18 7 D1
<< end >>
