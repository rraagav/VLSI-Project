magic
tech scmos
timestamp 1700492045
<< nwell >>
rect 323 49 383 73
rect 250 1 310 25
rect 424 -19 484 5
rect 492 -19 520 5
rect 338 -60 398 -36
<< ntransistor >>
rect 335 12 339 20
rect 356 12 360 20
rect 262 -36 266 -28
rect 283 -36 287 -28
rect 436 -56 440 -48
rect 457 -56 461 -48
rect 504 -50 508 -42
rect 350 -97 354 -89
rect 371 -97 375 -89
<< ptransistor >>
rect 335 57 339 65
rect 356 57 360 65
rect 262 9 266 17
rect 283 9 287 17
rect 436 -11 440 -3
rect 457 -11 461 -3
rect 504 -11 508 -3
rect 350 -52 354 -44
rect 371 -52 375 -44
<< ndiffusion >>
rect 329 18 335 20
rect 329 14 330 18
rect 334 14 335 18
rect 329 12 335 14
rect 339 12 356 20
rect 360 18 377 20
rect 360 14 363 18
rect 367 14 377 18
rect 360 12 377 14
rect 256 -30 262 -28
rect 256 -34 257 -30
rect 261 -34 262 -30
rect 256 -36 262 -34
rect 266 -36 283 -28
rect 287 -30 304 -28
rect 287 -34 290 -30
rect 294 -34 304 -30
rect 287 -36 304 -34
rect 498 -44 504 -42
rect 498 -48 499 -44
rect 503 -48 504 -44
rect 430 -50 436 -48
rect 430 -54 431 -50
rect 435 -54 436 -50
rect 430 -56 436 -54
rect 440 -56 457 -48
rect 461 -50 478 -48
rect 498 -50 504 -48
rect 508 -44 514 -42
rect 508 -48 509 -44
rect 513 -48 514 -44
rect 508 -50 514 -48
rect 461 -54 464 -50
rect 468 -54 478 -50
rect 461 -56 478 -54
rect 344 -91 350 -89
rect 344 -95 345 -91
rect 349 -95 350 -91
rect 344 -97 350 -95
rect 354 -97 371 -89
rect 375 -91 392 -89
rect 375 -95 378 -91
rect 382 -95 392 -91
rect 375 -97 392 -95
<< pdiffusion >>
rect 329 63 335 65
rect 329 59 330 63
rect 334 59 335 63
rect 329 57 335 59
rect 339 63 356 65
rect 339 59 340 63
rect 344 59 356 63
rect 339 57 356 59
rect 360 63 377 65
rect 360 59 363 63
rect 367 59 377 63
rect 360 57 377 59
rect 256 15 262 17
rect 256 11 257 15
rect 261 11 262 15
rect 256 9 262 11
rect 266 15 283 17
rect 266 11 267 15
rect 271 11 283 15
rect 266 9 283 11
rect 287 15 304 17
rect 287 11 290 15
rect 294 11 304 15
rect 287 9 304 11
rect 430 -5 436 -3
rect 430 -9 431 -5
rect 435 -9 436 -5
rect 430 -11 436 -9
rect 440 -5 457 -3
rect 440 -9 441 -5
rect 445 -9 457 -5
rect 440 -11 457 -9
rect 461 -5 478 -3
rect 461 -9 464 -5
rect 468 -9 478 -5
rect 461 -11 478 -9
rect 498 -5 504 -3
rect 498 -9 499 -5
rect 503 -9 504 -5
rect 498 -11 504 -9
rect 508 -5 514 -3
rect 508 -9 509 -5
rect 513 -9 514 -5
rect 508 -11 514 -9
rect 344 -46 350 -44
rect 344 -50 345 -46
rect 349 -50 350 -46
rect 344 -52 350 -50
rect 354 -46 371 -44
rect 354 -50 355 -46
rect 359 -50 371 -46
rect 354 -52 371 -50
rect 375 -46 392 -44
rect 375 -50 378 -46
rect 382 -50 392 -46
rect 375 -52 392 -50
<< ndcontact >>
rect 330 14 334 18
rect 363 14 367 18
rect 257 -34 261 -30
rect 290 -34 294 -30
rect 499 -48 503 -44
rect 431 -54 435 -50
rect 509 -48 513 -44
rect 464 -54 468 -50
rect 345 -95 349 -91
rect 378 -95 382 -91
<< pdcontact >>
rect 330 59 334 63
rect 340 59 344 63
rect 363 59 367 63
rect 257 11 261 15
rect 267 11 271 15
rect 290 11 294 15
rect 431 -9 435 -5
rect 441 -9 445 -5
rect 464 -9 468 -5
rect 499 -9 503 -5
rect 509 -9 513 -5
rect 345 -50 349 -46
rect 355 -50 359 -46
rect 378 -50 382 -46
<< polysilicon >>
rect 335 65 339 68
rect 356 65 360 68
rect 335 20 339 57
rect 356 20 360 57
rect 262 17 266 20
rect 283 17 287 20
rect 335 9 339 12
rect 262 -28 266 9
rect 283 -28 287 9
rect 356 5 360 12
rect 436 -3 440 0
rect 457 -3 461 0
rect 504 -3 508 0
rect 262 -39 266 -36
rect 283 -44 287 -36
rect 350 -44 354 -41
rect 371 -44 375 -41
rect 436 -48 440 -11
rect 457 -48 461 -11
rect 504 -42 508 -11
rect 350 -89 354 -52
rect 371 -89 375 -52
rect 504 -53 508 -50
rect 436 -59 440 -56
rect 457 -64 461 -56
rect 350 -100 354 -97
rect 371 -105 375 -97
<< polycontact >>
rect 331 38 335 42
rect 258 -10 262 -6
rect 352 4 356 8
rect 432 -30 436 -26
rect 279 -44 283 -40
rect 500 -34 504 -30
rect 346 -71 350 -67
rect 453 -64 457 -60
rect 367 -105 371 -101
<< metal1 >>
rect 299 81 468 85
rect 238 65 311 69
rect 238 -6 242 65
rect 307 42 311 65
rect 330 63 334 81
rect 363 63 367 81
rect 307 38 331 42
rect 340 38 344 59
rect 340 34 408 38
rect 257 30 294 34
rect 257 15 261 30
rect 290 15 294 30
rect 363 18 367 34
rect 234 -10 258 -6
rect 267 -10 271 11
rect 348 -10 352 8
rect 267 -14 352 -10
rect 290 -30 294 -14
rect 275 -67 279 -40
rect 267 -71 279 -67
rect 320 -67 324 -14
rect 345 -28 386 -24
rect 404 -26 408 34
rect 431 -5 435 81
rect 464 17 468 81
rect 464 13 503 17
rect 464 -5 468 13
rect 499 -5 503 13
rect 345 -46 349 -28
rect 378 -46 382 -28
rect 404 -30 432 -26
rect 441 -30 445 -9
rect 509 -30 513 -9
rect 441 -34 500 -30
rect 509 -34 521 -30
rect 464 -50 468 -34
rect 509 -44 513 -34
rect 320 -71 346 -67
rect 355 -71 359 -50
rect 499 -58 503 -48
rect 449 -71 453 -60
rect 492 -62 503 -58
rect 275 -120 279 -71
rect 355 -75 453 -71
rect 378 -91 382 -75
rect 363 -120 367 -101
rect 275 -124 367 -120
<< m2contact >>
rect 294 81 299 86
rect 289 34 294 39
rect 329 9 334 14
rect 256 -39 261 -34
rect 386 -28 391 -23
rect 426 15 431 20
rect 430 -59 435 -54
rect 492 -67 497 -62
rect 344 -100 349 -95
<< metal2 >>
rect 290 39 294 85
rect 391 15 426 19
rect 257 -48 261 -39
rect 330 -48 334 9
rect 391 -28 395 15
rect 250 -52 334 -48
rect 330 -109 334 -52
rect 431 -79 435 -59
rect 492 -79 496 -67
rect 431 -83 496 -79
rect 345 -109 349 -100
rect 431 -109 435 -83
rect 330 -113 435 -109
<< labels >>
rlabel metal1 268 -70 270 -69 1 VB
rlabel metal1 235 -8 237 -7 3 VA
rlabel metal2 251 -51 254 -49 1 GND
rlabel metal1 258 31 263 33 1 VDD
rlabel metal1 517 -33 520 -32 7 Vout
<< end >>
