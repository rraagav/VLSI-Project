magic
tech scmos
timestamp 1700504172
<< nwell >>
rect 21 0 81 24
rect 87 0 115 24
rect 21 -93 81 -69
rect 87 -93 115 -69
rect 21 -185 81 -161
rect 87 -185 115 -161
rect 21 -278 81 -254
rect 87 -278 115 -254
<< ntransistor >>
rect 33 -37 37 -29
rect 54 -37 58 -29
rect 99 -37 103 -29
rect 33 -130 37 -122
rect 54 -130 58 -122
rect 99 -130 103 -122
rect 33 -222 37 -214
rect 54 -222 58 -214
rect 99 -222 103 -214
rect 33 -315 37 -307
rect 54 -315 58 -307
rect 99 -315 103 -307
<< ptransistor >>
rect 33 8 37 16
rect 54 8 58 16
rect 99 8 103 16
rect 33 -85 37 -77
rect 54 -85 58 -77
rect 99 -85 103 -77
rect 33 -177 37 -169
rect 54 -177 58 -169
rect 99 -177 103 -169
rect 33 -270 37 -262
rect 54 -270 58 -262
rect 99 -270 103 -262
<< ndiffusion >>
rect 27 -31 33 -29
rect 27 -35 28 -31
rect 32 -35 33 -31
rect 27 -37 33 -35
rect 37 -37 54 -29
rect 58 -31 75 -29
rect 58 -35 61 -31
rect 65 -35 75 -31
rect 58 -37 75 -35
rect 93 -31 99 -29
rect 93 -35 94 -31
rect 98 -35 99 -31
rect 93 -37 99 -35
rect 103 -31 109 -29
rect 103 -35 104 -31
rect 108 -35 109 -31
rect 103 -37 109 -35
rect 27 -124 33 -122
rect 27 -128 28 -124
rect 32 -128 33 -124
rect 27 -130 33 -128
rect 37 -130 54 -122
rect 58 -124 75 -122
rect 58 -128 61 -124
rect 65 -128 75 -124
rect 58 -130 75 -128
rect 93 -124 99 -122
rect 93 -128 94 -124
rect 98 -128 99 -124
rect 93 -130 99 -128
rect 103 -124 109 -122
rect 103 -128 104 -124
rect 108 -128 109 -124
rect 103 -130 109 -128
rect 27 -216 33 -214
rect 27 -220 28 -216
rect 32 -220 33 -216
rect 27 -222 33 -220
rect 37 -222 54 -214
rect 58 -216 75 -214
rect 58 -220 61 -216
rect 65 -220 75 -216
rect 58 -222 75 -220
rect 93 -216 99 -214
rect 93 -220 94 -216
rect 98 -220 99 -216
rect 93 -222 99 -220
rect 103 -216 109 -214
rect 103 -220 104 -216
rect 108 -220 109 -216
rect 103 -222 109 -220
rect 27 -309 33 -307
rect 27 -313 28 -309
rect 32 -313 33 -309
rect 27 -315 33 -313
rect 37 -315 54 -307
rect 58 -309 75 -307
rect 58 -313 61 -309
rect 65 -313 75 -309
rect 58 -315 75 -313
rect 93 -309 99 -307
rect 93 -313 94 -309
rect 98 -313 99 -309
rect 93 -315 99 -313
rect 103 -309 109 -307
rect 103 -313 104 -309
rect 108 -313 109 -309
rect 103 -315 109 -313
<< pdiffusion >>
rect 27 14 33 16
rect 27 10 28 14
rect 32 10 33 14
rect 27 8 33 10
rect 37 14 54 16
rect 37 10 38 14
rect 42 10 54 14
rect 37 8 54 10
rect 58 14 75 16
rect 58 10 61 14
rect 65 10 75 14
rect 58 8 75 10
rect 93 14 99 16
rect 93 10 94 14
rect 98 10 99 14
rect 93 8 99 10
rect 103 14 109 16
rect 103 10 104 14
rect 108 10 109 14
rect 103 8 109 10
rect 27 -79 33 -77
rect 27 -83 28 -79
rect 32 -83 33 -79
rect 27 -85 33 -83
rect 37 -79 54 -77
rect 37 -83 38 -79
rect 42 -83 54 -79
rect 37 -85 54 -83
rect 58 -79 75 -77
rect 58 -83 61 -79
rect 65 -83 75 -79
rect 58 -85 75 -83
rect 93 -79 99 -77
rect 93 -83 94 -79
rect 98 -83 99 -79
rect 93 -85 99 -83
rect 103 -79 109 -77
rect 103 -83 104 -79
rect 108 -83 109 -79
rect 103 -85 109 -83
rect 27 -171 33 -169
rect 27 -175 28 -171
rect 32 -175 33 -171
rect 27 -177 33 -175
rect 37 -171 54 -169
rect 37 -175 38 -171
rect 42 -175 54 -171
rect 37 -177 54 -175
rect 58 -171 75 -169
rect 58 -175 61 -171
rect 65 -175 75 -171
rect 58 -177 75 -175
rect 93 -171 99 -169
rect 93 -175 94 -171
rect 98 -175 99 -171
rect 93 -177 99 -175
rect 103 -171 109 -169
rect 103 -175 104 -171
rect 108 -175 109 -171
rect 103 -177 109 -175
rect 27 -264 33 -262
rect 27 -268 28 -264
rect 32 -268 33 -264
rect 27 -270 33 -268
rect 37 -264 54 -262
rect 37 -268 38 -264
rect 42 -268 54 -264
rect 37 -270 54 -268
rect 58 -264 75 -262
rect 58 -268 61 -264
rect 65 -268 75 -264
rect 58 -270 75 -268
rect 93 -264 99 -262
rect 93 -268 94 -264
rect 98 -268 99 -264
rect 93 -270 99 -268
rect 103 -264 109 -262
rect 103 -268 104 -264
rect 108 -268 109 -264
rect 103 -270 109 -268
<< ndcontact >>
rect 28 -35 32 -31
rect 61 -35 65 -31
rect 94 -35 98 -31
rect 104 -35 108 -31
rect 28 -128 32 -124
rect 61 -128 65 -124
rect 94 -128 98 -124
rect 104 -128 108 -124
rect 28 -220 32 -216
rect 61 -220 65 -216
rect 94 -220 98 -216
rect 104 -220 108 -216
rect 28 -313 32 -309
rect 61 -313 65 -309
rect 94 -313 98 -309
rect 104 -313 108 -309
<< pdcontact >>
rect 28 10 32 14
rect 38 10 42 14
rect 61 10 65 14
rect 94 10 98 14
rect 104 10 108 14
rect 28 -83 32 -79
rect 38 -83 42 -79
rect 61 -83 65 -79
rect 94 -83 98 -79
rect 104 -83 108 -79
rect 28 -175 32 -171
rect 38 -175 42 -171
rect 61 -175 65 -171
rect 94 -175 98 -171
rect 104 -175 108 -171
rect 28 -268 32 -264
rect 38 -268 42 -264
rect 61 -268 65 -264
rect 94 -268 98 -264
rect 104 -268 108 -264
<< polysilicon >>
rect 33 16 37 19
rect 54 16 58 19
rect 99 16 103 19
rect 33 -29 37 8
rect 54 -29 58 8
rect 99 -29 103 8
rect 33 -40 37 -37
rect 54 -40 58 -37
rect 99 -40 103 -37
rect 33 -77 37 -74
rect 54 -77 58 -74
rect 99 -77 103 -74
rect 33 -122 37 -85
rect 54 -122 58 -85
rect 99 -122 103 -85
rect 33 -133 37 -130
rect 54 -133 58 -130
rect 99 -133 103 -130
rect 33 -169 37 -166
rect 54 -169 58 -166
rect 99 -169 103 -166
rect 33 -214 37 -177
rect 54 -214 58 -177
rect 99 -214 103 -177
rect 33 -225 37 -222
rect 54 -225 58 -222
rect 99 -225 103 -222
rect 33 -262 37 -259
rect 54 -262 58 -259
rect 99 -262 103 -259
rect 33 -307 37 -270
rect 54 -307 58 -270
rect 99 -307 103 -270
rect 33 -318 37 -315
rect 54 -318 58 -315
rect 99 -318 103 -315
<< polycontact >>
rect 29 -11 33 -7
rect 50 -23 54 -19
rect 95 -15 99 -11
rect 29 -104 33 -100
rect 50 -116 54 -112
rect 95 -108 99 -104
rect 29 -196 33 -192
rect 50 -208 54 -204
rect 95 -200 99 -196
rect 29 -289 33 -285
rect 50 -301 54 -297
rect 95 -293 99 -289
<< metal1 >>
rect 28 32 135 36
rect 28 14 32 32
rect 61 14 65 32
rect 94 14 98 32
rect 17 -11 29 -7
rect 38 -11 42 10
rect 38 -15 95 -11
rect 17 -23 50 -19
rect 61 -31 65 -15
rect 104 -16 108 10
rect 104 -20 115 -16
rect 104 -31 108 -20
rect 28 -45 32 -35
rect 94 -45 98 -35
rect 28 -49 98 -45
rect 131 -57 135 32
rect 28 -61 135 -57
rect 28 -79 32 -61
rect 61 -79 65 -61
rect 94 -79 98 -61
rect 17 -104 29 -100
rect 38 -104 42 -83
rect 38 -108 95 -104
rect 17 -116 50 -112
rect 61 -124 65 -108
rect 104 -109 108 -83
rect 104 -113 115 -109
rect 104 -124 108 -113
rect 28 -138 32 -128
rect 94 -138 98 -128
rect 28 -142 98 -138
rect 131 -149 135 -61
rect 28 -153 135 -149
rect 28 -171 32 -153
rect 61 -171 65 -153
rect 94 -171 98 -153
rect 17 -196 29 -192
rect 38 -196 42 -175
rect 38 -200 95 -196
rect 17 -208 50 -204
rect 61 -216 65 -200
rect 104 -201 108 -175
rect 104 -205 115 -201
rect 104 -216 108 -205
rect 28 -230 32 -220
rect 94 -230 98 -220
rect 28 -234 98 -230
rect 131 -242 135 -153
rect 28 -246 135 -242
rect 28 -264 32 -246
rect 61 -264 65 -246
rect 94 -264 98 -246
rect 17 -289 29 -285
rect 38 -289 42 -268
rect 38 -293 95 -289
rect 17 -301 50 -297
rect 61 -309 65 -293
rect 104 -294 108 -268
rect 104 -298 115 -294
rect 104 -309 108 -298
rect 28 -323 32 -313
rect 94 -323 98 -313
rect 28 -327 98 -323
<< m2contact >>
rect 98 -49 103 -44
rect 98 -142 103 -137
rect 98 -234 103 -229
rect 98 -327 103 -322
<< metal2 >>
rect 103 -49 127 -45
rect 123 -138 127 -49
rect 103 -142 127 -138
rect 123 -230 127 -142
rect 103 -234 127 -230
rect 123 -323 127 -234
rect 103 -327 127 -323
<< labels >>
rlabel metal1 18 -10 20 -9 1 A0
rlabel metal1 18 -22 20 -21 1 B0
rlabel metal1 18 -103 20 -102 3 A1
rlabel metal1 18 -115 20 -114 3 B1
rlabel metal1 111 -19 113 -18 1 Ans0
rlabel metal1 31 34 34 35 5 VDD
rlabel metal1 111 -112 113 -111 1 Ans1
rlabel metal1 32 -48 35 -47 1 GND
rlabel metal1 18 -196 21 -194 3 A2
rlabel metal1 18 -207 21 -205 3 B2
rlabel metal1 18 -288 21 -286 3 A3
rlabel metal1 18 -300 20 -299 3 B3
rlabel metal1 111 -204 113 -203 1 Ans2
rlabel metal1 111 -297 113 -296 1 Ans3
<< end >>
