* SPICE3 file created from 3and.ext - technology: scmos
.include TSMC_180nm.txt

.param SUPPLY = 1.8
.param LAMBDA = 0.18u
.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}
.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd VDD gnd 'Supply'

* Vin_VA VA gnd PULSE(0 1.8 0ns 200ps 200ps 199ns 400ns)
* Vin_VB VB gnd PULSE(0 1.8 0ns 200ps 200ps 399ns 800ns)
* Vin_VC VC gnd PULSE(0 1.8 0ns 200ps 200ps 599ns 1000ns)

Vin_VC VC gnd DC(1.8)
Vin_VB VB gnd DC(1.8)
Vin_VA VA gnd DC(1.8)

.option scale=0.09u

M1000 a_14_8# VC a_43_n44# Gnd CMOSN w=8 l=4
+  ad=144 pd=52 as=160 ps=56
M1001 Vout a_14_8# VDD w_99_0# CMOSP w=8 l=4
+  ad=48 pd=28 as=256 ps=112
M1002 Vout a_14_8# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=96 ps=56
M1003 a_14_n44# VA GND Gnd CMOSN w=8 l=4
+  ad=200 pd=66 as=0 ps=0
M1004 a_14_8# VC VDD w_n2_0# CMOSP w=8 l=4
+  ad=344 pd=118 as=0 ps=0
M1005 a_43_n44# VB a_14_n44# Gnd CMOSN w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1006 a_14_8# VA VDD w_n2_0# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1007 VDD VB a_14_8# w_n2_0# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
C0 w_n2_0# VA 0.11fF
C1 VDD Vout 0.03fF
C2 VA a_14_8# 0.03fF
C3 w_99_0# VDD 0.03fF
C4 VB VC 0.49fF
C5 w_n2_0# VC 0.11fF
C6 Vout GND 0.03fF
C7 VC GND 0.03fF
C8 a_14_8# Vout 0.03fF
C9 VC a_14_8# 0.10fF
C10 w_n2_0# VDD 0.05fF
C11 VA VC 0.10fF
C12 w_99_0# a_14_8# 0.11fF
C13 w_n2_0# VB 0.11fF
C14 a_14_8# VDD 0.03fF
C15 w_99_0# Vout 0.03fF
C16 VB a_14_8# 0.35fF
C17 VA VB 0.10fF
C18 w_n2_0# a_14_8# 0.05fF
C19 Vout Gnd 0.14fF
C20 a_14_8# Gnd 0.76fF
C21 VC Gnd 0.52fF
C22 VB Gnd 0.45fF
C23 VA Gnd 0.37fF
C24 w_99_0# Gnd 0.67fF
C25 w_n2_0# Gnd 2.24fF

.tran 1n 1600n
.control
run
plot v(VA) v(VB)+2 v(VC)+4 v(Vout)+6
.end
.endc