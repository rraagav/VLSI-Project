magic
tech scmos
timestamp 1700488508
<< nwell >>
rect -2 0 58 24
<< ntransistor >>
rect 10 -40 14 -32
rect 31 -40 35 -32
<< ptransistor >>
rect 10 8 14 16
rect 31 8 35 16
<< ndiffusion >>
rect 4 -34 10 -32
rect 4 -38 5 -34
rect 9 -38 10 -34
rect 4 -40 10 -38
rect 14 -34 31 -32
rect 14 -38 15 -34
rect 19 -38 31 -34
rect 14 -40 31 -38
rect 35 -34 52 -32
rect 35 -38 38 -34
rect 42 -38 52 -34
rect 35 -40 52 -38
<< pdiffusion >>
rect 4 14 10 16
rect 4 10 5 14
rect 9 10 10 14
rect 4 8 10 10
rect 14 8 31 16
rect 35 14 52 16
rect 35 10 40 14
rect 44 10 52 14
rect 35 8 52 10
<< ndcontact >>
rect 5 -38 9 -34
rect 15 -38 19 -34
rect 38 -38 42 -34
<< pdcontact >>
rect 5 10 9 14
rect 40 10 44 14
<< polysilicon >>
rect 10 16 14 19
rect 31 16 35 19
rect 10 -32 14 8
rect 31 -32 35 8
rect 10 -43 14 -40
rect 31 -43 35 -40
<< polycontact >>
rect 6 -12 10 -8
rect 27 -20 31 -16
<< metal1 >>
rect -2 32 25 36
rect 5 14 9 32
rect 2 -12 6 -8
rect 2 -20 27 -16
rect 40 -24 44 10
rect 15 -28 58 -24
rect 15 -34 19 -28
rect 5 -50 9 -38
rect 38 -50 42 -38
rect -2 -54 42 -50
<< labels >>
rlabel metal1 2 34 4 35 4 VDD
rlabel metal1 3 -11 5 -10 1 VA
rlabel metal1 2 -53 4 -52 2 GND
rlabel metal1 51 -27 54 -26 1 Vout
rlabel metal1 3 -19 5 -18 1 VB
<< end >>
