* SPICE3 file created from or.ext - technology: scmos
.include TSMC_180nm.txt

.param SUPPLY = 1.8
.param LAMBDA = 0.18u
.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}
.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd VDD gnd 'Supply'

Vin_A VA gnd DC(1.8)
Vin_B VB gnd DC(1.8)

* Vin_VA VA gnd PULSE(0 1.8 0ns 100ps 100ps 199ns 400ns)
* Vin_VB VB gnd PULSE(0 1.8 0ns 100ps 100ps 399ns 800ns)

.option scale=0.09u

M1000 Vout a_88_n46# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=232 ps=106
M1001 a_88_2# VA VDD w_72_n6# CMOSP w=8 l=4
+  ad=136 pd=50 as=96 ps=56
M1002 a_88_n46# VB a_88_2# w_72_n6# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1003 Vout a_88_n46# VDD w_140_n6# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1004 a_88_n46# VA GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1005 GND VB a_88_n46# Gnd CMOSN w=8 l=4
+  ad=0 pd=0 as=0 ps=0
C0 w_72_n6# VB 0.11fF
C1 a_88_n46# Vout 0.03fF
C2 w_140_n6# Vout 0.03fF
C3 w_72_n6# VDD 0.03fF
C4 VA VB 0.19fF
C5 w_140_n6# a_88_n46# 0.11fF
C6 w_72_n6# VA 0.11fF
C7 VB a_88_n46# 0.27fF
C8 w_72_n6# a_88_n46# 0.03fF
C9 Vout GND 0.03fF
C10 a_88_n46# GND 0.08fF
C11 VDD Vout 0.03fF
C12 w_140_n6# VDD 0.03fF
C13 GND Gnd 0.35fF
C14 Vout Gnd 0.11fF
C15 VDD Gnd 0.31fF
C16 a_88_n46# Gnd 0.59fF
C17 VB Gnd 0.40fF
C18 VA Gnd 0.34fF
C19 w_140_n6# Gnd 0.55fF
C20 w_72_n6# Gnd 1.45fF

.tran 1n 800n
.control
run
plot v(Vout)+4 v(VB)+2 v(VA)
.end
.endc