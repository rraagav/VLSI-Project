magic
tech scmos
timestamp 1700521080
<< nwell >>
rect 71 44 131 68
rect 560 44 620 68
rect 944 44 1004 68
rect 1359 20 1419 44
rect -2 -4 58 20
rect 172 -24 232 0
rect 487 -4 547 20
rect 298 -28 326 -4
rect 661 -24 721 0
rect 871 -4 931 20
rect 734 -28 762 -4
rect 1079 -24 1139 0
rect 1152 -28 1180 -4
rect 1286 -28 1346 -4
rect 86 -65 146 -41
rect 575 -65 635 -41
rect 959 -65 1019 -41
rect 1460 -48 1520 -24
rect 1528 -48 1556 -24
rect 1374 -89 1434 -65
rect 391 -314 488 -290
rect 499 -314 527 -290
rect 807 -314 904 -290
rect 915 -314 943 -290
rect 1257 -314 1354 -290
rect 1365 -314 1393 -290
rect 313 -367 341 -343
rect 729 -367 757 -343
rect 1173 -367 1201 -343
rect 24 -391 52 -367
rect 111 -399 171 -375
rect 177 -399 205 -375
rect 313 -459 341 -435
rect 409 -451 506 -427
rect 517 -451 545 -427
rect 22 -484 50 -460
rect 722 -487 750 -463
rect 825 -479 922 -455
rect 933 -479 961 -455
rect 1172 -459 1200 -435
rect 1275 -451 1372 -427
rect 1383 -451 1411 -427
rect 112 -515 172 -491
rect 178 -515 206 -491
rect 1014 -497 1074 -473
rect 1080 -497 1108 -473
rect 1495 -492 1611 -468
rect 1619 -492 1647 -468
rect 605 -536 665 -512
rect 671 -536 699 -512
rect 93 -693 216 -669
rect 224 -693 252 -669
rect 363 -693 486 -669
rect 494 -693 522 -669
<< ntransistor >>
rect 83 7 87 15
rect 104 7 108 15
rect 572 7 576 15
rect 593 7 597 15
rect 10 -41 14 -33
rect 31 -41 35 -33
rect 956 7 960 15
rect 977 7 981 15
rect 499 -41 503 -33
rect 520 -41 524 -33
rect 184 -61 188 -53
rect 205 -61 209 -53
rect 310 -59 314 -51
rect 883 -41 887 -33
rect 904 -41 908 -33
rect 673 -61 677 -53
rect 694 -61 698 -53
rect 746 -59 750 -51
rect 1371 -17 1375 -9
rect 1392 -17 1396 -9
rect 1091 -61 1095 -53
rect 1112 -61 1116 -53
rect 1164 -59 1168 -51
rect 1298 -65 1302 -57
rect 1319 -65 1323 -57
rect 98 -102 102 -94
rect 119 -102 123 -94
rect 587 -102 591 -94
rect 608 -102 612 -94
rect 971 -102 975 -94
rect 992 -102 996 -94
rect 1472 -85 1476 -77
rect 1493 -85 1497 -77
rect 1540 -79 1544 -71
rect 1386 -126 1390 -118
rect 1407 -126 1411 -118
rect 36 -422 40 -414
rect 403 -380 407 -372
rect 436 -380 440 -372
rect 460 -380 464 -372
rect 511 -380 515 -372
rect 819 -380 823 -372
rect 852 -380 856 -372
rect 876 -380 880 -372
rect 927 -380 931 -372
rect 1269 -380 1273 -372
rect 1302 -380 1306 -372
rect 1326 -380 1330 -372
rect 1377 -380 1381 -372
rect 325 -404 329 -396
rect 741 -404 745 -396
rect 1185 -404 1189 -396
rect 123 -436 127 -428
rect 144 -436 148 -428
rect 189 -436 193 -428
rect 325 -496 329 -488
rect 34 -515 38 -507
rect 421 -517 425 -509
rect 454 -517 458 -509
rect 478 -517 482 -509
rect 529 -517 533 -509
rect 734 -524 738 -516
rect 124 -552 128 -544
rect 145 -552 149 -544
rect 190 -552 194 -544
rect 1184 -496 1188 -488
rect 1287 -517 1291 -509
rect 1320 -517 1324 -509
rect 1344 -517 1348 -509
rect 1395 -517 1399 -509
rect 1026 -534 1030 -526
rect 1047 -534 1051 -526
rect 1092 -534 1096 -526
rect 837 -545 841 -537
rect 870 -545 874 -537
rect 894 -545 898 -537
rect 945 -545 949 -537
rect 1507 -546 1511 -538
rect 1536 -546 1540 -538
rect 1560 -546 1564 -538
rect 1584 -546 1588 -538
rect 1631 -546 1635 -538
rect 617 -573 621 -565
rect 638 -573 642 -565
rect 683 -573 687 -565
rect 105 -753 109 -745
rect 126 -753 130 -745
rect 147 -753 151 -745
rect 168 -753 172 -745
rect 236 -753 240 -745
rect 375 -756 379 -748
rect 396 -756 400 -748
rect 417 -756 421 -748
rect 438 -756 442 -748
rect 506 -756 510 -748
<< ptransistor >>
rect 83 52 87 60
rect 104 52 108 60
rect 572 52 576 60
rect 593 52 597 60
rect 956 52 960 60
rect 977 52 981 60
rect 1371 28 1375 36
rect 1392 28 1396 36
rect 10 4 14 12
rect 31 4 35 12
rect 499 4 503 12
rect 520 4 524 12
rect 184 -16 188 -8
rect 205 -16 209 -8
rect 98 -57 102 -49
rect 119 -57 123 -49
rect 310 -20 314 -12
rect 883 4 887 12
rect 904 4 908 12
rect 673 -16 677 -8
rect 694 -16 698 -8
rect 587 -57 591 -49
rect 608 -57 612 -49
rect 746 -20 750 -12
rect 1091 -16 1095 -8
rect 1112 -16 1116 -8
rect 971 -57 975 -49
rect 992 -57 996 -49
rect 1164 -20 1168 -12
rect 1298 -20 1302 -12
rect 1319 -20 1323 -12
rect 1472 -40 1476 -32
rect 1493 -40 1497 -32
rect 1540 -40 1544 -32
rect 1386 -81 1390 -73
rect 1407 -81 1411 -73
rect 403 -306 407 -298
rect 436 -306 440 -298
rect 460 -306 464 -298
rect 511 -306 515 -298
rect 819 -306 823 -298
rect 852 -306 856 -298
rect 876 -306 880 -298
rect 927 -306 931 -298
rect 1269 -306 1273 -298
rect 1302 -306 1306 -298
rect 1326 -306 1330 -298
rect 1377 -306 1381 -298
rect 325 -359 329 -351
rect 36 -383 40 -375
rect 123 -391 127 -383
rect 144 -391 148 -383
rect 189 -391 193 -383
rect 741 -359 745 -351
rect 1185 -359 1189 -351
rect 421 -443 425 -435
rect 454 -443 458 -435
rect 478 -443 482 -435
rect 529 -443 533 -435
rect 325 -451 329 -443
rect 34 -476 38 -468
rect 124 -507 128 -499
rect 145 -507 149 -499
rect 190 -507 194 -499
rect 1287 -443 1291 -435
rect 1320 -443 1324 -435
rect 1344 -443 1348 -435
rect 1395 -443 1399 -435
rect 1184 -451 1188 -443
rect 837 -471 841 -463
rect 870 -471 874 -463
rect 894 -471 898 -463
rect 945 -471 949 -463
rect 734 -479 738 -471
rect 617 -528 621 -520
rect 638 -528 642 -520
rect 683 -528 687 -520
rect 1026 -489 1030 -481
rect 1047 -489 1051 -481
rect 1092 -489 1096 -481
rect 1507 -484 1511 -476
rect 1536 -484 1540 -476
rect 1560 -484 1564 -476
rect 1584 -484 1588 -476
rect 1631 -484 1635 -476
rect 105 -685 109 -677
rect 126 -685 130 -677
rect 147 -685 151 -677
rect 168 -685 172 -677
rect 236 -685 240 -677
rect 375 -685 379 -677
rect 396 -685 400 -677
rect 417 -685 421 -677
rect 438 -685 442 -677
rect 506 -685 510 -677
<< ndiffusion >>
rect 77 13 83 15
rect 77 9 78 13
rect 82 9 83 13
rect 77 7 83 9
rect 87 7 104 15
rect 108 13 125 15
rect 108 9 111 13
rect 115 9 125 13
rect 566 13 572 15
rect 108 7 125 9
rect 566 9 567 13
rect 571 9 572 13
rect 566 7 572 9
rect 576 7 593 15
rect 597 13 614 15
rect 597 9 600 13
rect 604 9 614 13
rect 950 13 956 15
rect 597 7 614 9
rect 4 -35 10 -33
rect 4 -39 5 -35
rect 9 -39 10 -35
rect 4 -41 10 -39
rect 14 -41 31 -33
rect 35 -35 52 -33
rect 35 -39 38 -35
rect 42 -39 52 -35
rect 35 -41 52 -39
rect 950 9 951 13
rect 955 9 956 13
rect 950 7 956 9
rect 960 7 977 15
rect 981 13 998 15
rect 981 9 984 13
rect 988 9 998 13
rect 981 7 998 9
rect 493 -35 499 -33
rect 493 -39 494 -35
rect 498 -39 499 -35
rect 493 -41 499 -39
rect 503 -41 520 -33
rect 524 -35 541 -33
rect 524 -39 527 -35
rect 531 -39 541 -35
rect 524 -41 541 -39
rect 304 -53 310 -51
rect 178 -55 184 -53
rect 178 -59 179 -55
rect 183 -59 184 -55
rect 178 -61 184 -59
rect 188 -61 205 -53
rect 209 -55 226 -53
rect 209 -59 212 -55
rect 216 -59 226 -55
rect 304 -57 305 -53
rect 309 -57 310 -53
rect 304 -59 310 -57
rect 314 -53 320 -51
rect 314 -57 315 -53
rect 319 -57 320 -53
rect 1365 -11 1371 -9
rect 877 -35 883 -33
rect 877 -39 878 -35
rect 882 -39 883 -35
rect 877 -41 883 -39
rect 887 -41 904 -33
rect 908 -35 925 -33
rect 908 -39 911 -35
rect 915 -39 925 -35
rect 908 -41 925 -39
rect 740 -53 746 -51
rect 667 -55 673 -53
rect 314 -59 320 -57
rect 209 -61 226 -59
rect 667 -59 668 -55
rect 672 -59 673 -55
rect 667 -61 673 -59
rect 677 -61 694 -53
rect 698 -55 715 -53
rect 698 -59 701 -55
rect 705 -59 715 -55
rect 740 -57 741 -53
rect 745 -57 746 -53
rect 740 -59 746 -57
rect 750 -53 756 -51
rect 750 -57 751 -53
rect 755 -57 756 -53
rect 1365 -15 1366 -11
rect 1370 -15 1371 -11
rect 1365 -17 1371 -15
rect 1375 -17 1392 -9
rect 1396 -11 1413 -9
rect 1396 -15 1399 -11
rect 1403 -15 1413 -11
rect 1396 -17 1413 -15
rect 1158 -53 1164 -51
rect 1085 -55 1091 -53
rect 750 -59 756 -57
rect 698 -61 715 -59
rect 1085 -59 1086 -55
rect 1090 -59 1091 -55
rect 1085 -61 1091 -59
rect 1095 -61 1112 -53
rect 1116 -55 1133 -53
rect 1116 -59 1119 -55
rect 1123 -59 1133 -55
rect 1158 -57 1159 -53
rect 1163 -57 1164 -53
rect 1158 -59 1164 -57
rect 1168 -53 1174 -51
rect 1168 -57 1169 -53
rect 1173 -57 1174 -53
rect 1168 -59 1174 -57
rect 1292 -59 1298 -57
rect 1116 -61 1133 -59
rect 1292 -63 1293 -59
rect 1297 -63 1298 -59
rect 1292 -65 1298 -63
rect 1302 -65 1319 -57
rect 1323 -59 1340 -57
rect 1323 -63 1326 -59
rect 1330 -63 1340 -59
rect 1323 -65 1340 -63
rect 1534 -73 1540 -71
rect 1534 -77 1535 -73
rect 1539 -77 1540 -73
rect 1466 -79 1472 -77
rect 92 -96 98 -94
rect 92 -100 93 -96
rect 97 -100 98 -96
rect 92 -102 98 -100
rect 102 -102 119 -94
rect 123 -96 140 -94
rect 123 -100 126 -96
rect 130 -100 140 -96
rect 123 -102 140 -100
rect 581 -96 587 -94
rect 581 -100 582 -96
rect 586 -100 587 -96
rect 581 -102 587 -100
rect 591 -102 608 -94
rect 612 -96 629 -94
rect 612 -100 615 -96
rect 619 -100 629 -96
rect 612 -102 629 -100
rect 965 -96 971 -94
rect 965 -100 966 -96
rect 970 -100 971 -96
rect 965 -102 971 -100
rect 975 -102 992 -94
rect 996 -96 1013 -94
rect 996 -100 999 -96
rect 1003 -100 1013 -96
rect 996 -102 1013 -100
rect -55 -115 -39 -107
rect 1466 -83 1467 -79
rect 1471 -83 1472 -79
rect 1466 -85 1472 -83
rect 1476 -85 1493 -77
rect 1497 -79 1514 -77
rect 1534 -79 1540 -77
rect 1544 -73 1550 -71
rect 1544 -77 1545 -73
rect 1549 -77 1550 -73
rect 1544 -79 1550 -77
rect 1497 -83 1500 -79
rect 1504 -83 1514 -79
rect 1497 -85 1514 -83
rect 1380 -120 1386 -118
rect 1380 -124 1381 -120
rect 1385 -124 1386 -120
rect 1380 -126 1386 -124
rect 1390 -126 1407 -118
rect 1411 -120 1428 -118
rect 1411 -124 1414 -120
rect 1418 -124 1428 -120
rect 1411 -126 1428 -124
rect -106 -215 -101 -207
rect -138 -232 -133 -224
rect -149 -257 -144 -249
rect 30 -416 36 -414
rect 30 -420 31 -416
rect 35 -420 36 -416
rect 30 -422 36 -420
rect 40 -416 46 -414
rect 40 -420 41 -416
rect 45 -420 46 -416
rect 40 -422 46 -420
rect 397 -374 403 -372
rect 397 -378 398 -374
rect 402 -378 403 -374
rect 397 -380 403 -378
rect 407 -380 436 -372
rect 440 -380 460 -372
rect 464 -374 482 -372
rect 464 -378 471 -374
rect 475 -378 482 -374
rect 464 -380 482 -378
rect 505 -374 511 -372
rect 505 -378 506 -374
rect 510 -378 511 -374
rect 505 -380 511 -378
rect 515 -374 521 -372
rect 515 -378 516 -374
rect 520 -378 521 -374
rect 515 -380 521 -378
rect 813 -374 819 -372
rect 813 -378 814 -374
rect 818 -378 819 -374
rect 813 -380 819 -378
rect 823 -380 852 -372
rect 856 -380 876 -372
rect 880 -374 898 -372
rect 880 -378 887 -374
rect 891 -378 898 -374
rect 880 -380 898 -378
rect 921 -374 927 -372
rect 921 -378 922 -374
rect 926 -378 927 -374
rect 921 -380 927 -378
rect 931 -374 937 -372
rect 931 -378 932 -374
rect 936 -378 937 -374
rect 931 -380 937 -378
rect 1263 -374 1269 -372
rect 1263 -378 1264 -374
rect 1268 -378 1269 -374
rect 1263 -380 1269 -378
rect 1273 -380 1302 -372
rect 1306 -380 1326 -372
rect 1330 -374 1348 -372
rect 1330 -378 1337 -374
rect 1341 -378 1348 -374
rect 1330 -380 1348 -378
rect 1371 -374 1377 -372
rect 1371 -378 1372 -374
rect 1376 -378 1377 -374
rect 1371 -380 1377 -378
rect 1381 -374 1387 -372
rect 1381 -378 1382 -374
rect 1386 -378 1387 -374
rect 1381 -380 1387 -378
rect 319 -398 325 -396
rect 319 -402 320 -398
rect 324 -402 325 -398
rect 319 -404 325 -402
rect 329 -398 335 -396
rect 329 -402 330 -398
rect 334 -402 335 -398
rect 329 -404 335 -402
rect 735 -398 741 -396
rect 735 -402 736 -398
rect 740 -402 741 -398
rect 735 -404 741 -402
rect 745 -398 751 -396
rect 745 -402 746 -398
rect 750 -402 751 -398
rect 745 -404 751 -402
rect 1179 -398 1185 -396
rect 1179 -402 1180 -398
rect 1184 -402 1185 -398
rect 1179 -404 1185 -402
rect 1189 -398 1195 -396
rect 1189 -402 1190 -398
rect 1194 -402 1195 -398
rect 1189 -404 1195 -402
rect 259 -419 264 -414
rect 1116 -419 1121 -414
rect 117 -430 123 -428
rect 117 -434 118 -430
rect 122 -434 123 -430
rect 117 -436 123 -434
rect 127 -436 144 -428
rect 148 -430 165 -428
rect 148 -434 151 -430
rect 155 -434 165 -430
rect 148 -436 165 -434
rect 183 -430 189 -428
rect 183 -434 184 -430
rect 188 -434 189 -430
rect 183 -436 189 -434
rect 193 -430 199 -428
rect 193 -434 194 -430
rect 198 -434 199 -430
rect 193 -436 199 -434
rect 319 -490 325 -488
rect 319 -494 320 -490
rect 324 -494 325 -490
rect 319 -496 325 -494
rect 329 -490 335 -488
rect 329 -494 330 -490
rect 334 -494 335 -490
rect 329 -496 335 -494
rect 28 -509 34 -507
rect 28 -513 29 -509
rect 33 -513 34 -509
rect 28 -515 34 -513
rect 38 -509 44 -507
rect 38 -513 39 -509
rect 43 -513 44 -509
rect 38 -515 44 -513
rect 100 -540 105 -535
rect 672 -447 677 -442
rect 415 -511 421 -509
rect 415 -515 416 -511
rect 420 -515 421 -511
rect 415 -517 421 -515
rect 425 -517 454 -509
rect 458 -517 478 -509
rect 482 -511 500 -509
rect 482 -515 489 -511
rect 493 -515 500 -511
rect 482 -517 500 -515
rect 523 -511 529 -509
rect 523 -515 524 -511
rect 528 -515 529 -511
rect 523 -517 529 -515
rect 533 -511 539 -509
rect 533 -515 534 -511
rect 538 -515 539 -511
rect 533 -517 539 -515
rect 728 -518 734 -516
rect 728 -522 729 -518
rect 733 -522 734 -518
rect 728 -524 734 -522
rect 738 -518 744 -516
rect 738 -522 739 -518
rect 743 -522 744 -518
rect 738 -524 744 -522
rect 118 -546 124 -544
rect 118 -550 119 -546
rect 123 -550 124 -546
rect 118 -552 124 -550
rect 128 -552 145 -544
rect 149 -546 166 -544
rect 149 -550 152 -546
rect 156 -550 166 -546
rect 149 -552 166 -550
rect 184 -546 190 -544
rect 184 -550 185 -546
rect 189 -550 190 -546
rect 184 -552 190 -550
rect 194 -546 200 -544
rect 194 -550 195 -546
rect 199 -550 200 -546
rect 194 -552 200 -550
rect 1178 -490 1184 -488
rect 1178 -494 1179 -490
rect 1183 -494 1184 -490
rect 1178 -496 1184 -494
rect 1188 -490 1194 -488
rect 1188 -494 1189 -490
rect 1193 -494 1194 -490
rect 1188 -496 1194 -494
rect 1281 -511 1287 -509
rect 1281 -515 1282 -511
rect 1286 -515 1287 -511
rect 1281 -517 1287 -515
rect 1291 -517 1320 -509
rect 1324 -517 1344 -509
rect 1348 -511 1366 -509
rect 1348 -515 1355 -511
rect 1359 -515 1366 -511
rect 1348 -517 1366 -515
rect 1389 -511 1395 -509
rect 1389 -515 1390 -511
rect 1394 -515 1395 -511
rect 1389 -517 1395 -515
rect 1399 -511 1405 -509
rect 1399 -515 1400 -511
rect 1404 -515 1405 -511
rect 1399 -517 1405 -515
rect 1020 -528 1026 -526
rect 1020 -532 1021 -528
rect 1025 -532 1026 -528
rect 1020 -534 1026 -532
rect 1030 -534 1047 -526
rect 1051 -528 1068 -526
rect 1051 -532 1054 -528
rect 1058 -532 1068 -528
rect 1051 -534 1068 -532
rect 1086 -528 1092 -526
rect 1086 -532 1087 -528
rect 1091 -532 1092 -528
rect 1086 -534 1092 -532
rect 1096 -528 1102 -526
rect 1096 -532 1097 -528
rect 1101 -532 1102 -528
rect 1096 -534 1102 -532
rect 831 -539 837 -537
rect 831 -543 832 -539
rect 836 -543 837 -539
rect 831 -545 837 -543
rect 841 -545 870 -537
rect 874 -545 894 -537
rect 898 -539 916 -537
rect 898 -543 905 -539
rect 909 -543 916 -539
rect 898 -545 916 -543
rect 939 -539 945 -537
rect 939 -543 940 -539
rect 944 -543 945 -539
rect 939 -545 945 -543
rect 949 -539 955 -537
rect 949 -543 950 -539
rect 954 -543 955 -539
rect 949 -545 955 -543
rect 1501 -540 1507 -538
rect 1501 -544 1502 -540
rect 1506 -544 1507 -540
rect 1501 -546 1507 -544
rect 1511 -546 1536 -538
rect 1540 -546 1560 -538
rect 1564 -546 1584 -538
rect 1588 -540 1605 -538
rect 1588 -544 1594 -540
rect 1598 -544 1605 -540
rect 1588 -546 1605 -544
rect 1625 -540 1631 -538
rect 1625 -544 1626 -540
rect 1630 -544 1631 -540
rect 1625 -546 1631 -544
rect 1635 -540 1641 -538
rect 1635 -544 1636 -540
rect 1640 -544 1641 -540
rect 1635 -546 1641 -544
rect 611 -567 617 -565
rect 611 -571 612 -567
rect 616 -571 617 -567
rect 611 -573 617 -571
rect 621 -573 638 -565
rect 642 -567 659 -565
rect 642 -571 645 -567
rect 649 -571 659 -567
rect 642 -573 659 -571
rect 677 -567 683 -565
rect 677 -571 678 -567
rect 682 -571 683 -567
rect 677 -573 683 -571
rect 687 -567 693 -565
rect 687 -571 688 -567
rect 692 -571 693 -567
rect 687 -573 693 -571
rect 99 -747 105 -745
rect 99 -751 100 -747
rect 104 -751 105 -747
rect 99 -753 105 -751
rect 109 -747 126 -745
rect 109 -751 110 -747
rect 114 -751 126 -747
rect 109 -753 126 -751
rect 130 -747 147 -745
rect 130 -751 133 -747
rect 137 -751 147 -747
rect 130 -753 147 -751
rect 151 -747 168 -745
rect 151 -751 157 -747
rect 161 -751 168 -747
rect 151 -753 168 -751
rect 172 -753 210 -745
rect 230 -747 236 -745
rect 230 -751 231 -747
rect 235 -751 236 -747
rect 230 -753 236 -751
rect 240 -747 246 -745
rect 240 -751 241 -747
rect 245 -751 246 -747
rect 240 -753 246 -751
rect 369 -750 375 -748
rect 369 -754 370 -750
rect 374 -754 375 -750
rect 369 -756 375 -754
rect 379 -750 396 -748
rect 379 -754 380 -750
rect 384 -754 396 -750
rect 379 -756 396 -754
rect 400 -750 417 -748
rect 400 -754 403 -750
rect 407 -754 417 -750
rect 400 -756 417 -754
rect 421 -750 438 -748
rect 421 -754 427 -750
rect 431 -754 438 -750
rect 421 -756 438 -754
rect 442 -756 480 -748
rect 500 -750 506 -748
rect 500 -754 501 -750
rect 505 -754 506 -750
rect 500 -756 506 -754
rect 510 -750 516 -748
rect 510 -754 511 -750
rect 515 -754 516 -750
rect 510 -756 516 -754
<< pdiffusion >>
rect 77 58 83 60
rect 77 54 78 58
rect 82 54 83 58
rect 77 52 83 54
rect 87 58 104 60
rect 87 54 88 58
rect 92 54 104 58
rect 87 52 104 54
rect 108 58 125 60
rect 108 54 111 58
rect 115 54 125 58
rect 108 52 125 54
rect 566 58 572 60
rect 566 54 567 58
rect 571 54 572 58
rect 566 52 572 54
rect 576 58 593 60
rect 576 54 577 58
rect 581 54 593 58
rect 576 52 593 54
rect 597 58 614 60
rect 597 54 600 58
rect 604 54 614 58
rect 597 52 614 54
rect 950 58 956 60
rect 950 54 951 58
rect 955 54 956 58
rect 950 52 956 54
rect 960 58 977 60
rect 960 54 961 58
rect 965 54 977 58
rect 960 52 977 54
rect 981 58 998 60
rect 981 54 984 58
rect 988 54 998 58
rect 981 52 998 54
rect 1365 34 1371 36
rect 1365 30 1366 34
rect 1370 30 1371 34
rect 1365 28 1371 30
rect 1375 34 1392 36
rect 1375 30 1376 34
rect 1380 30 1392 34
rect 1375 28 1392 30
rect 1396 34 1413 36
rect 1396 30 1399 34
rect 1403 30 1413 34
rect 1396 28 1413 30
rect 4 10 10 12
rect 4 6 5 10
rect 9 6 10 10
rect 4 4 10 6
rect 14 10 31 12
rect 14 6 15 10
rect 19 6 31 10
rect 14 4 31 6
rect 35 10 52 12
rect 35 6 38 10
rect 42 6 52 10
rect 493 10 499 12
rect 35 4 52 6
rect 493 6 494 10
rect 498 6 499 10
rect 493 4 499 6
rect 503 10 520 12
rect 503 6 504 10
rect 508 6 520 10
rect 503 4 520 6
rect 524 10 541 12
rect 524 6 527 10
rect 531 6 541 10
rect 877 10 883 12
rect 524 4 541 6
rect 178 -10 184 -8
rect 178 -14 179 -10
rect 183 -14 184 -10
rect 178 -16 184 -14
rect 188 -10 205 -8
rect 188 -14 189 -10
rect 193 -14 205 -10
rect 188 -16 205 -14
rect 209 -10 226 -8
rect 209 -14 212 -10
rect 216 -14 226 -10
rect 209 -16 226 -14
rect 304 -14 310 -12
rect 92 -51 98 -49
rect 92 -55 93 -51
rect 97 -55 98 -51
rect 92 -57 98 -55
rect 102 -51 119 -49
rect 102 -55 103 -51
rect 107 -55 119 -51
rect 102 -57 119 -55
rect 123 -51 140 -49
rect 123 -55 126 -51
rect 130 -55 140 -51
rect 304 -18 305 -14
rect 309 -18 310 -14
rect 304 -20 310 -18
rect 314 -14 320 -12
rect 314 -18 315 -14
rect 319 -18 320 -14
rect 314 -20 320 -18
rect 877 6 878 10
rect 882 6 883 10
rect 877 4 883 6
rect 887 10 904 12
rect 887 6 888 10
rect 892 6 904 10
rect 887 4 904 6
rect 908 10 925 12
rect 908 6 911 10
rect 915 6 925 10
rect 908 4 925 6
rect 667 -10 673 -8
rect 667 -14 668 -10
rect 672 -14 673 -10
rect 667 -16 673 -14
rect 677 -10 694 -8
rect 677 -14 678 -10
rect 682 -14 694 -10
rect 677 -16 694 -14
rect 698 -10 715 -8
rect 698 -14 701 -10
rect 705 -14 715 -10
rect 698 -16 715 -14
rect 740 -14 746 -12
rect 581 -51 587 -49
rect 123 -57 140 -55
rect 581 -55 582 -51
rect 586 -55 587 -51
rect 581 -57 587 -55
rect 591 -51 608 -49
rect 591 -55 592 -51
rect 596 -55 608 -51
rect 591 -57 608 -55
rect 612 -51 629 -49
rect 612 -55 615 -51
rect 619 -55 629 -51
rect 740 -18 741 -14
rect 745 -18 746 -14
rect 740 -20 746 -18
rect 750 -14 756 -12
rect 750 -18 751 -14
rect 755 -18 756 -14
rect 750 -20 756 -18
rect 1085 -10 1091 -8
rect 1085 -14 1086 -10
rect 1090 -14 1091 -10
rect 1085 -16 1091 -14
rect 1095 -10 1112 -8
rect 1095 -14 1096 -10
rect 1100 -14 1112 -10
rect 1095 -16 1112 -14
rect 1116 -10 1133 -8
rect 1116 -14 1119 -10
rect 1123 -14 1133 -10
rect 1116 -16 1133 -14
rect 1158 -14 1164 -12
rect 965 -51 971 -49
rect 612 -57 629 -55
rect 965 -55 966 -51
rect 970 -55 971 -51
rect 965 -57 971 -55
rect 975 -51 992 -49
rect 975 -55 976 -51
rect 980 -55 992 -51
rect 975 -57 992 -55
rect 996 -51 1013 -49
rect 996 -55 999 -51
rect 1003 -55 1013 -51
rect 1158 -18 1159 -14
rect 1163 -18 1164 -14
rect 1158 -20 1164 -18
rect 1168 -14 1174 -12
rect 1168 -18 1169 -14
rect 1173 -18 1174 -14
rect 1168 -20 1174 -18
rect 1292 -14 1298 -12
rect 1292 -18 1293 -14
rect 1297 -18 1298 -14
rect 1292 -20 1298 -18
rect 1302 -14 1319 -12
rect 1302 -18 1303 -14
rect 1307 -18 1319 -14
rect 1302 -20 1319 -18
rect 1323 -14 1340 -12
rect 1323 -18 1326 -14
rect 1330 -18 1340 -14
rect 1323 -20 1340 -18
rect 996 -57 1013 -55
rect 1466 -34 1472 -32
rect 1466 -38 1467 -34
rect 1471 -38 1472 -34
rect 1466 -40 1472 -38
rect 1476 -34 1493 -32
rect 1476 -38 1477 -34
rect 1481 -38 1493 -34
rect 1476 -40 1493 -38
rect 1497 -34 1514 -32
rect 1497 -38 1500 -34
rect 1504 -38 1514 -34
rect 1497 -40 1514 -38
rect 1534 -34 1540 -32
rect 1534 -38 1535 -34
rect 1539 -38 1540 -34
rect 1534 -40 1540 -38
rect 1544 -34 1550 -32
rect 1544 -38 1545 -34
rect 1549 -38 1550 -34
rect 1544 -40 1550 -38
rect 1380 -75 1386 -73
rect 1380 -79 1381 -75
rect 1385 -79 1386 -75
rect 1380 -81 1386 -79
rect 1390 -75 1407 -73
rect 1390 -79 1391 -75
rect 1395 -79 1407 -75
rect 1390 -81 1407 -79
rect 1411 -75 1428 -73
rect 1411 -79 1414 -75
rect 1418 -79 1428 -75
rect 1411 -81 1428 -79
rect 397 -300 403 -298
rect 397 -304 398 -300
rect 402 -304 403 -300
rect 397 -306 403 -304
rect 407 -300 436 -298
rect 407 -304 412 -300
rect 416 -304 436 -300
rect 407 -306 436 -304
rect 440 -300 460 -298
rect 440 -304 453 -300
rect 457 -304 460 -300
rect 440 -306 460 -304
rect 464 -300 482 -298
rect 464 -304 471 -300
rect 475 -304 482 -300
rect 464 -306 482 -304
rect 505 -300 511 -298
rect 505 -304 506 -300
rect 510 -304 511 -300
rect 505 -306 511 -304
rect 515 -300 521 -298
rect 515 -304 516 -300
rect 520 -304 521 -300
rect 515 -306 521 -304
rect 813 -300 819 -298
rect 813 -304 814 -300
rect 818 -304 819 -300
rect 813 -306 819 -304
rect 823 -300 852 -298
rect 823 -304 828 -300
rect 832 -304 852 -300
rect 823 -306 852 -304
rect 856 -300 876 -298
rect 856 -304 869 -300
rect 873 -304 876 -300
rect 856 -306 876 -304
rect 880 -300 898 -298
rect 880 -304 887 -300
rect 891 -304 898 -300
rect 880 -306 898 -304
rect 921 -300 927 -298
rect 921 -304 922 -300
rect 926 -304 927 -300
rect 921 -306 927 -304
rect 931 -300 937 -298
rect 931 -304 932 -300
rect 936 -304 937 -300
rect 931 -306 937 -304
rect 1263 -300 1269 -298
rect 1263 -304 1264 -300
rect 1268 -304 1269 -300
rect 1263 -306 1269 -304
rect 1273 -300 1302 -298
rect 1273 -304 1278 -300
rect 1282 -304 1302 -300
rect 1273 -306 1302 -304
rect 1306 -300 1326 -298
rect 1306 -304 1319 -300
rect 1323 -304 1326 -300
rect 1306 -306 1326 -304
rect 1330 -300 1348 -298
rect 1330 -304 1337 -300
rect 1341 -304 1348 -300
rect 1330 -306 1348 -304
rect 1371 -300 1377 -298
rect 1371 -304 1372 -300
rect 1376 -304 1377 -300
rect 1371 -306 1377 -304
rect 1381 -300 1387 -298
rect 1381 -304 1382 -300
rect 1386 -304 1387 -300
rect 1381 -306 1387 -304
rect 319 -353 325 -351
rect 319 -357 320 -353
rect 324 -357 325 -353
rect 319 -359 325 -357
rect 329 -353 335 -351
rect 329 -357 330 -353
rect 334 -357 335 -353
rect 329 -359 335 -357
rect 30 -377 36 -375
rect 30 -381 31 -377
rect 35 -381 36 -377
rect 30 -383 36 -381
rect 40 -377 46 -375
rect 40 -381 41 -377
rect 45 -381 46 -377
rect 40 -383 46 -381
rect 117 -385 123 -383
rect 117 -389 118 -385
rect 122 -389 123 -385
rect 117 -391 123 -389
rect 127 -385 144 -383
rect 127 -389 128 -385
rect 132 -389 144 -385
rect 127 -391 144 -389
rect 148 -385 165 -383
rect 148 -389 151 -385
rect 155 -389 165 -385
rect 148 -391 165 -389
rect 183 -385 189 -383
rect 183 -389 184 -385
rect 188 -389 189 -385
rect 183 -391 189 -389
rect 193 -385 199 -383
rect 193 -389 194 -385
rect 198 -389 199 -385
rect 193 -391 199 -389
rect 735 -353 741 -351
rect 735 -357 736 -353
rect 740 -357 741 -353
rect 735 -359 741 -357
rect 745 -353 751 -351
rect 745 -357 746 -353
rect 750 -357 751 -353
rect 745 -359 751 -357
rect 1179 -353 1185 -351
rect 1179 -357 1180 -353
rect 1184 -357 1185 -353
rect 1179 -359 1185 -357
rect 1189 -353 1195 -351
rect 1189 -357 1190 -353
rect 1194 -357 1195 -353
rect 1189 -359 1195 -357
rect 415 -437 421 -435
rect 415 -441 416 -437
rect 420 -441 421 -437
rect 415 -443 421 -441
rect 425 -437 454 -435
rect 425 -441 430 -437
rect 434 -441 454 -437
rect 425 -443 454 -441
rect 458 -437 478 -435
rect 458 -441 471 -437
rect 475 -441 478 -437
rect 458 -443 478 -441
rect 482 -437 500 -435
rect 482 -441 489 -437
rect 493 -441 500 -437
rect 482 -443 500 -441
rect 523 -437 529 -435
rect 523 -441 524 -437
rect 528 -441 529 -437
rect 523 -443 529 -441
rect 533 -437 539 -435
rect 533 -441 534 -437
rect 538 -441 539 -437
rect 1281 -437 1287 -435
rect 533 -443 539 -441
rect 319 -445 325 -443
rect 319 -449 320 -445
rect 324 -449 325 -445
rect 319 -451 325 -449
rect 329 -445 335 -443
rect 329 -449 330 -445
rect 334 -449 335 -445
rect 329 -451 335 -449
rect 28 -470 34 -468
rect 28 -474 29 -470
rect 33 -474 34 -470
rect 28 -476 34 -474
rect 38 -470 44 -468
rect 38 -474 39 -470
rect 43 -474 44 -470
rect 38 -476 44 -474
rect 118 -501 124 -499
rect 118 -505 119 -501
rect 123 -505 124 -501
rect 118 -507 124 -505
rect 128 -501 145 -499
rect 128 -505 129 -501
rect 133 -505 145 -501
rect 128 -507 145 -505
rect 149 -501 166 -499
rect 149 -505 152 -501
rect 156 -505 166 -501
rect 149 -507 166 -505
rect 184 -501 190 -499
rect 184 -505 185 -501
rect 189 -505 190 -501
rect 184 -507 190 -505
rect 194 -501 200 -499
rect 194 -505 195 -501
rect 199 -505 200 -501
rect 194 -507 200 -505
rect 1281 -441 1282 -437
rect 1286 -441 1287 -437
rect 1281 -443 1287 -441
rect 1291 -437 1320 -435
rect 1291 -441 1296 -437
rect 1300 -441 1320 -437
rect 1291 -443 1320 -441
rect 1324 -437 1344 -435
rect 1324 -441 1337 -437
rect 1341 -441 1344 -437
rect 1324 -443 1344 -441
rect 1348 -437 1366 -435
rect 1348 -441 1355 -437
rect 1359 -441 1366 -437
rect 1348 -443 1366 -441
rect 1389 -437 1395 -435
rect 1389 -441 1390 -437
rect 1394 -441 1395 -437
rect 1389 -443 1395 -441
rect 1399 -437 1405 -435
rect 1399 -441 1400 -437
rect 1404 -441 1405 -437
rect 1399 -443 1405 -441
rect 1178 -445 1184 -443
rect 1178 -449 1179 -445
rect 1183 -449 1184 -445
rect 1178 -451 1184 -449
rect 1188 -445 1194 -443
rect 1188 -449 1189 -445
rect 1193 -449 1194 -445
rect 1188 -451 1194 -449
rect 831 -465 837 -463
rect 831 -469 832 -465
rect 836 -469 837 -465
rect 831 -471 837 -469
rect 841 -465 870 -463
rect 841 -469 846 -465
rect 850 -469 870 -465
rect 841 -471 870 -469
rect 874 -465 894 -463
rect 874 -469 887 -465
rect 891 -469 894 -465
rect 874 -471 894 -469
rect 898 -465 916 -463
rect 898 -469 905 -465
rect 909 -469 916 -465
rect 898 -471 916 -469
rect 939 -465 945 -463
rect 939 -469 940 -465
rect 944 -469 945 -465
rect 939 -471 945 -469
rect 949 -465 955 -463
rect 949 -469 950 -465
rect 954 -469 955 -465
rect 949 -471 955 -469
rect 728 -473 734 -471
rect 728 -477 729 -473
rect 733 -477 734 -473
rect 728 -479 734 -477
rect 738 -473 744 -471
rect 738 -477 739 -473
rect 743 -477 744 -473
rect 738 -479 744 -477
rect 611 -522 617 -520
rect 611 -526 612 -522
rect 616 -526 617 -522
rect 611 -528 617 -526
rect 621 -522 638 -520
rect 621 -526 622 -522
rect 626 -526 638 -522
rect 621 -528 638 -526
rect 642 -522 659 -520
rect 642 -526 645 -522
rect 649 -526 659 -522
rect 642 -528 659 -526
rect 677 -522 683 -520
rect 677 -526 678 -522
rect 682 -526 683 -522
rect 677 -528 683 -526
rect 687 -522 693 -520
rect 687 -526 688 -522
rect 692 -526 693 -522
rect 687 -528 693 -526
rect 1020 -483 1026 -481
rect 1020 -487 1021 -483
rect 1025 -487 1026 -483
rect 1020 -489 1026 -487
rect 1030 -483 1047 -481
rect 1030 -487 1031 -483
rect 1035 -487 1047 -483
rect 1030 -489 1047 -487
rect 1051 -483 1068 -481
rect 1051 -487 1054 -483
rect 1058 -487 1068 -483
rect 1051 -489 1068 -487
rect 1086 -483 1092 -481
rect 1086 -487 1087 -483
rect 1091 -487 1092 -483
rect 1086 -489 1092 -487
rect 1096 -483 1102 -481
rect 1096 -487 1097 -483
rect 1101 -487 1102 -483
rect 1096 -489 1102 -487
rect 1501 -478 1507 -476
rect 1501 -482 1502 -478
rect 1506 -482 1507 -478
rect 1501 -484 1507 -482
rect 1511 -478 1536 -476
rect 1511 -482 1512 -478
rect 1516 -482 1536 -478
rect 1511 -484 1536 -482
rect 1540 -478 1560 -476
rect 1540 -482 1553 -478
rect 1557 -482 1560 -478
rect 1540 -484 1560 -482
rect 1564 -478 1584 -476
rect 1564 -482 1573 -478
rect 1577 -482 1584 -478
rect 1564 -484 1584 -482
rect 1588 -478 1605 -476
rect 1588 -482 1594 -478
rect 1598 -482 1605 -478
rect 1588 -484 1605 -482
rect 1625 -478 1631 -476
rect 1625 -482 1626 -478
rect 1630 -482 1631 -478
rect 1625 -484 1631 -482
rect 1635 -478 1641 -476
rect 1635 -482 1636 -478
rect 1640 -482 1641 -478
rect 1635 -484 1641 -482
rect 99 -679 105 -677
rect 99 -683 100 -679
rect 104 -683 105 -679
rect 99 -685 105 -683
rect 109 -685 126 -677
rect 130 -685 147 -677
rect 151 -685 168 -677
rect 172 -679 210 -677
rect 172 -683 184 -679
rect 188 -683 210 -679
rect 172 -685 210 -683
rect 230 -679 236 -677
rect 230 -683 231 -679
rect 235 -683 236 -679
rect 230 -685 236 -683
rect 240 -679 246 -677
rect 240 -683 241 -679
rect 245 -683 246 -679
rect 240 -685 246 -683
rect 369 -679 375 -677
rect 369 -683 370 -679
rect 374 -683 375 -679
rect 369 -685 375 -683
rect 379 -685 396 -677
rect 400 -685 417 -677
rect 421 -685 438 -677
rect 442 -679 480 -677
rect 442 -683 454 -679
rect 458 -683 480 -679
rect 442 -685 480 -683
rect 500 -679 506 -677
rect 500 -683 501 -679
rect 505 -683 506 -679
rect 500 -685 506 -683
rect 510 -679 516 -677
rect 510 -683 511 -679
rect 515 -683 516 -679
rect 510 -685 516 -683
<< ndcontact >>
rect 78 9 82 13
rect 111 9 115 13
rect 567 9 571 13
rect 600 9 604 13
rect 5 -39 9 -35
rect 38 -39 42 -35
rect 951 9 955 13
rect 984 9 988 13
rect 494 -39 498 -35
rect 527 -39 531 -35
rect 179 -59 183 -55
rect 212 -59 216 -55
rect 305 -57 309 -53
rect 315 -57 319 -53
rect 878 -39 882 -35
rect 911 -39 915 -35
rect 668 -59 672 -55
rect 701 -59 705 -55
rect 741 -57 745 -53
rect 751 -57 755 -53
rect 1366 -15 1370 -11
rect 1399 -15 1403 -11
rect 1086 -59 1090 -55
rect 1119 -59 1123 -55
rect 1159 -57 1163 -53
rect 1169 -57 1173 -53
rect 1293 -63 1297 -59
rect 1326 -63 1330 -59
rect 1535 -77 1539 -73
rect 93 -100 97 -96
rect 126 -100 130 -96
rect 582 -100 586 -96
rect 615 -100 619 -96
rect 966 -100 970 -96
rect 999 -100 1003 -96
rect 1467 -83 1471 -79
rect 1545 -77 1549 -73
rect 1500 -83 1504 -79
rect 1381 -124 1385 -120
rect 1414 -124 1418 -120
rect 31 -420 35 -416
rect 41 -420 45 -416
rect 398 -378 402 -374
rect 471 -378 475 -374
rect 506 -378 510 -374
rect 516 -378 520 -374
rect 814 -378 818 -374
rect 887 -378 891 -374
rect 922 -378 926 -374
rect 932 -378 936 -374
rect 1264 -378 1268 -374
rect 1337 -378 1341 -374
rect 1372 -378 1376 -374
rect 1382 -378 1386 -374
rect 320 -402 324 -398
rect 330 -402 334 -398
rect 736 -402 740 -398
rect 746 -402 750 -398
rect 1180 -402 1184 -398
rect 1190 -402 1194 -398
rect 118 -434 122 -430
rect 151 -434 155 -430
rect 184 -434 188 -430
rect 194 -434 198 -430
rect 320 -494 324 -490
rect 330 -494 334 -490
rect 29 -513 33 -509
rect 39 -513 43 -509
rect 416 -515 420 -511
rect 489 -515 493 -511
rect 524 -515 528 -511
rect 534 -515 538 -511
rect 729 -522 733 -518
rect 739 -522 743 -518
rect 119 -550 123 -546
rect 152 -550 156 -546
rect 185 -550 189 -546
rect 195 -550 199 -546
rect 1179 -494 1183 -490
rect 1189 -494 1193 -490
rect 1282 -515 1286 -511
rect 1355 -515 1359 -511
rect 1390 -515 1394 -511
rect 1400 -515 1404 -511
rect 1021 -532 1025 -528
rect 1054 -532 1058 -528
rect 1087 -532 1091 -528
rect 1097 -532 1101 -528
rect 832 -543 836 -539
rect 905 -543 909 -539
rect 940 -543 944 -539
rect 950 -543 954 -539
rect 1502 -544 1506 -540
rect 1594 -544 1598 -540
rect 1626 -544 1630 -540
rect 1636 -544 1640 -540
rect 612 -571 616 -567
rect 645 -571 649 -567
rect 678 -571 682 -567
rect 688 -571 692 -567
rect 100 -751 104 -747
rect 110 -751 114 -747
rect 133 -751 137 -747
rect 157 -751 161 -747
rect 231 -751 235 -747
rect 241 -751 245 -747
rect 370 -754 374 -750
rect 380 -754 384 -750
rect 403 -754 407 -750
rect 427 -754 431 -750
rect 501 -754 505 -750
rect 511 -754 515 -750
<< pdcontact >>
rect 78 54 82 58
rect 88 54 92 58
rect 111 54 115 58
rect 567 54 571 58
rect 577 54 581 58
rect 600 54 604 58
rect 951 54 955 58
rect 961 54 965 58
rect 984 54 988 58
rect 1366 30 1370 34
rect 1376 30 1380 34
rect 1399 30 1403 34
rect 5 6 9 10
rect 15 6 19 10
rect 38 6 42 10
rect 494 6 498 10
rect 504 6 508 10
rect 527 6 531 10
rect 179 -14 183 -10
rect 189 -14 193 -10
rect 212 -14 216 -10
rect 93 -55 97 -51
rect 103 -55 107 -51
rect 126 -55 130 -51
rect 305 -18 309 -14
rect 315 -18 319 -14
rect 878 6 882 10
rect 888 6 892 10
rect 911 6 915 10
rect 668 -14 672 -10
rect 678 -14 682 -10
rect 701 -14 705 -10
rect 582 -55 586 -51
rect 592 -55 596 -51
rect 615 -55 619 -51
rect 741 -18 745 -14
rect 751 -18 755 -14
rect 1086 -14 1090 -10
rect 1096 -14 1100 -10
rect 1119 -14 1123 -10
rect 966 -55 970 -51
rect 976 -55 980 -51
rect 999 -55 1003 -51
rect 1159 -18 1163 -14
rect 1169 -18 1173 -14
rect 1293 -18 1297 -14
rect 1303 -18 1307 -14
rect 1326 -18 1330 -14
rect 1467 -38 1471 -34
rect 1477 -38 1481 -34
rect 1500 -38 1504 -34
rect 1535 -38 1539 -34
rect 1545 -38 1549 -34
rect 1381 -79 1385 -75
rect 1391 -79 1395 -75
rect 1414 -79 1418 -75
rect 398 -304 402 -300
rect 412 -304 416 -300
rect 453 -304 457 -300
rect 471 -304 475 -300
rect 506 -304 510 -300
rect 516 -304 520 -300
rect 814 -304 818 -300
rect 828 -304 832 -300
rect 869 -304 873 -300
rect 887 -304 891 -300
rect 922 -304 926 -300
rect 932 -304 936 -300
rect 1264 -304 1268 -300
rect 1278 -304 1282 -300
rect 1319 -304 1323 -300
rect 1337 -304 1341 -300
rect 1372 -304 1376 -300
rect 1382 -304 1386 -300
rect 320 -357 324 -353
rect 330 -357 334 -353
rect 31 -381 35 -377
rect 41 -381 45 -377
rect 118 -389 122 -385
rect 128 -389 132 -385
rect 151 -389 155 -385
rect 184 -389 188 -385
rect 194 -389 198 -385
rect 736 -357 740 -353
rect 746 -357 750 -353
rect 1180 -357 1184 -353
rect 1190 -357 1194 -353
rect 416 -441 420 -437
rect 430 -441 434 -437
rect 471 -441 475 -437
rect 489 -441 493 -437
rect 524 -441 528 -437
rect 534 -441 538 -437
rect 320 -449 324 -445
rect 330 -449 334 -445
rect 29 -474 33 -470
rect 39 -474 43 -470
rect 119 -505 123 -501
rect 129 -505 133 -501
rect 152 -505 156 -501
rect 185 -505 189 -501
rect 195 -505 199 -501
rect 1282 -441 1286 -437
rect 1296 -441 1300 -437
rect 1337 -441 1341 -437
rect 1355 -441 1359 -437
rect 1390 -441 1394 -437
rect 1400 -441 1404 -437
rect 1179 -449 1183 -445
rect 1189 -449 1193 -445
rect 832 -469 836 -465
rect 846 -469 850 -465
rect 887 -469 891 -465
rect 905 -469 909 -465
rect 940 -469 944 -465
rect 950 -469 954 -465
rect 729 -477 733 -473
rect 739 -477 743 -473
rect 612 -526 616 -522
rect 622 -526 626 -522
rect 645 -526 649 -522
rect 678 -526 682 -522
rect 688 -526 692 -522
rect 1021 -487 1025 -483
rect 1031 -487 1035 -483
rect 1054 -487 1058 -483
rect 1087 -487 1091 -483
rect 1097 -487 1101 -483
rect 1502 -482 1506 -478
rect 1512 -482 1516 -478
rect 1553 -482 1557 -478
rect 1573 -482 1577 -478
rect 1594 -482 1598 -478
rect 1626 -482 1630 -478
rect 1636 -482 1640 -478
rect 100 -683 104 -679
rect 184 -683 188 -679
rect 231 -683 235 -679
rect 241 -683 245 -679
rect 370 -683 374 -679
rect 454 -683 458 -679
rect 501 -683 505 -679
rect 511 -683 515 -679
<< polysilicon >>
rect 83 60 87 63
rect 104 60 108 63
rect 572 60 576 63
rect 593 60 597 63
rect 956 60 960 63
rect 977 60 981 63
rect 83 15 87 52
rect 104 15 108 52
rect 572 15 576 52
rect 593 15 597 52
rect 956 15 960 52
rect 977 15 981 52
rect 1371 36 1375 39
rect 1392 36 1396 39
rect 10 12 14 15
rect 31 12 35 15
rect 499 12 503 15
rect 520 12 524 15
rect 83 4 87 7
rect 10 -33 14 4
rect 31 -33 35 4
rect 104 0 108 7
rect 883 12 887 15
rect 904 12 908 15
rect 572 4 576 7
rect 184 -8 188 -5
rect 205 -8 209 -5
rect 310 -12 314 -9
rect 10 -44 14 -41
rect 31 -49 35 -41
rect 98 -49 102 -46
rect 119 -49 123 -46
rect 184 -53 188 -16
rect 205 -53 209 -16
rect 310 -51 314 -20
rect 499 -33 503 4
rect 520 -33 524 4
rect 593 0 597 7
rect 956 4 960 7
rect 673 -8 677 -5
rect 694 -8 698 -5
rect 746 -12 750 -9
rect 499 -44 503 -41
rect 520 -49 524 -41
rect 587 -49 591 -46
rect 608 -49 612 -46
rect 98 -94 102 -57
rect 119 -94 123 -57
rect 673 -53 677 -16
rect 694 -53 698 -16
rect 746 -51 750 -20
rect 883 -33 887 4
rect 904 -33 908 4
rect 977 0 981 7
rect 1091 -8 1095 -5
rect 1112 -8 1116 -5
rect 1371 -9 1375 28
rect 1392 -9 1396 28
rect 1164 -12 1168 -9
rect 1298 -12 1302 -9
rect 1319 -12 1323 -9
rect 883 -44 887 -41
rect 904 -49 908 -41
rect 971 -49 975 -46
rect 992 -49 996 -46
rect 184 -64 188 -61
rect 205 -69 209 -61
rect 310 -62 314 -59
rect 587 -94 591 -57
rect 608 -94 612 -57
rect 1091 -53 1095 -16
rect 1112 -53 1116 -16
rect 1371 -20 1375 -17
rect 1164 -51 1168 -20
rect 673 -64 677 -61
rect 694 -69 698 -61
rect 746 -62 750 -59
rect 971 -94 975 -57
rect 992 -94 996 -57
rect 1298 -57 1302 -20
rect 1319 -57 1323 -20
rect 1392 -24 1396 -17
rect 1472 -32 1476 -29
rect 1493 -32 1497 -29
rect 1540 -32 1544 -29
rect 1091 -64 1095 -61
rect 1112 -69 1116 -61
rect 1164 -62 1168 -59
rect 1298 -68 1302 -65
rect 1319 -73 1323 -65
rect 1386 -73 1390 -70
rect 1407 -73 1411 -70
rect 1472 -77 1476 -40
rect 1493 -77 1497 -40
rect 1540 -71 1544 -40
rect 98 -105 102 -102
rect 119 -110 123 -102
rect 587 -105 591 -102
rect 608 -110 612 -102
rect 971 -105 975 -102
rect 992 -110 996 -102
rect 1386 -118 1390 -81
rect 1407 -118 1411 -81
rect 1540 -82 1544 -79
rect 1472 -88 1476 -85
rect 1493 -93 1497 -85
rect 1386 -129 1390 -126
rect 1407 -134 1411 -126
rect 403 -298 407 -295
rect 436 -298 440 -295
rect 460 -298 464 -295
rect 511 -298 515 -295
rect 819 -298 823 -295
rect 852 -298 856 -295
rect 876 -298 880 -295
rect 927 -298 931 -295
rect 1269 -298 1273 -295
rect 1302 -298 1306 -295
rect 1326 -298 1330 -295
rect 1377 -298 1381 -295
rect 325 -351 329 -348
rect 36 -375 40 -372
rect 123 -383 127 -380
rect 144 -383 148 -380
rect 189 -383 193 -380
rect 36 -414 40 -383
rect 36 -425 40 -422
rect 123 -428 127 -391
rect 144 -428 148 -391
rect 189 -428 193 -391
rect 325 -396 329 -359
rect 403 -372 407 -306
rect 436 -372 440 -306
rect 460 -372 464 -306
rect 511 -372 515 -306
rect 741 -351 745 -348
rect 403 -383 407 -380
rect 436 -383 440 -380
rect 460 -383 464 -380
rect 511 -383 515 -380
rect 741 -396 745 -359
rect 819 -372 823 -306
rect 852 -372 856 -306
rect 876 -372 880 -306
rect 927 -372 931 -306
rect 1185 -351 1189 -348
rect 819 -383 823 -380
rect 852 -383 856 -380
rect 876 -383 880 -380
rect 927 -383 931 -380
rect 1185 -396 1189 -359
rect 1269 -372 1273 -306
rect 1302 -372 1306 -306
rect 1326 -372 1330 -306
rect 1377 -372 1381 -306
rect 1269 -383 1273 -380
rect 1302 -383 1306 -380
rect 1326 -383 1330 -380
rect 1377 -383 1381 -380
rect 325 -407 329 -404
rect 741 -407 745 -404
rect 1185 -407 1189 -404
rect 421 -435 425 -432
rect 454 -435 458 -432
rect 478 -435 482 -432
rect 529 -435 533 -432
rect 1287 -435 1291 -432
rect 1320 -435 1324 -432
rect 1344 -435 1348 -432
rect 1395 -435 1399 -432
rect 123 -439 127 -436
rect 144 -444 148 -436
rect 189 -439 193 -436
rect 325 -443 329 -440
rect 34 -468 38 -465
rect 34 -507 38 -476
rect 325 -488 329 -451
rect 124 -499 128 -496
rect 145 -499 149 -496
rect 190 -499 194 -496
rect 325 -499 329 -496
rect 34 -518 38 -515
rect 124 -544 128 -507
rect 145 -544 149 -507
rect 190 -544 194 -507
rect 421 -509 425 -443
rect 454 -509 458 -443
rect 478 -509 482 -443
rect 529 -509 533 -443
rect 1184 -443 1188 -440
rect 837 -463 841 -460
rect 870 -463 874 -460
rect 894 -463 898 -460
rect 945 -463 949 -460
rect 734 -471 738 -468
rect 734 -516 738 -479
rect 421 -520 425 -517
rect 454 -520 458 -517
rect 478 -520 482 -517
rect 529 -520 533 -517
rect 617 -520 621 -517
rect 638 -520 642 -517
rect 683 -520 687 -517
rect 734 -527 738 -524
rect 124 -555 128 -552
rect 145 -560 149 -552
rect 190 -555 194 -552
rect 617 -565 621 -528
rect 638 -565 642 -528
rect 683 -565 687 -528
rect 837 -537 841 -471
rect 870 -537 874 -471
rect 894 -537 898 -471
rect 945 -537 949 -471
rect 1026 -481 1030 -478
rect 1047 -481 1051 -478
rect 1092 -481 1096 -478
rect 1184 -488 1188 -451
rect 1026 -526 1030 -489
rect 1047 -526 1051 -489
rect 1092 -526 1096 -489
rect 1184 -499 1188 -496
rect 1287 -509 1291 -443
rect 1320 -509 1324 -443
rect 1344 -509 1348 -443
rect 1395 -509 1399 -443
rect 1507 -476 1511 -473
rect 1536 -476 1540 -473
rect 1560 -476 1564 -473
rect 1584 -476 1588 -473
rect 1631 -476 1635 -473
rect 1287 -520 1291 -517
rect 1320 -520 1324 -517
rect 1344 -520 1348 -517
rect 1395 -520 1399 -517
rect 1026 -537 1030 -534
rect 1047 -537 1051 -534
rect 1092 -537 1096 -534
rect 1507 -538 1511 -484
rect 1536 -538 1540 -484
rect 1560 -538 1564 -484
rect 1584 -538 1588 -484
rect 1631 -538 1635 -484
rect 837 -548 841 -545
rect 870 -548 874 -545
rect 894 -548 898 -545
rect 945 -548 949 -545
rect 1507 -549 1511 -546
rect 1536 -549 1540 -546
rect 1560 -549 1564 -546
rect 1584 -549 1588 -546
rect 1631 -549 1635 -546
rect 617 -576 621 -573
rect 638 -576 642 -573
rect 683 -576 687 -573
rect 105 -677 109 -674
rect 126 -677 130 -674
rect 147 -677 151 -674
rect 168 -677 172 -674
rect 236 -677 240 -674
rect 375 -677 379 -674
rect 396 -677 400 -674
rect 417 -677 421 -674
rect 438 -677 442 -674
rect 506 -677 510 -674
rect 105 -745 109 -685
rect 126 -745 130 -685
rect 147 -745 151 -685
rect 168 -745 172 -685
rect 236 -745 240 -685
rect 375 -748 379 -685
rect 396 -748 400 -685
rect 417 -748 421 -685
rect 438 -748 442 -685
rect 506 -748 510 -685
rect 105 -756 109 -753
rect 126 -756 130 -753
rect 147 -756 151 -753
rect 168 -756 172 -753
rect 236 -756 240 -753
rect 375 -759 379 -756
rect 396 -759 400 -756
rect 417 -759 421 -756
rect 438 -759 442 -756
rect 506 -759 510 -756
<< polycontact >>
rect 79 33 83 37
rect 568 33 572 37
rect 952 33 956 37
rect 6 -15 10 -11
rect 100 -1 104 3
rect 180 -35 184 -31
rect 27 -49 31 -45
rect 495 -19 499 -11
rect 306 -39 310 -35
rect 589 -1 593 3
rect 1367 9 1371 13
rect 669 -35 673 -31
rect 516 -49 520 -45
rect 94 -76 98 -72
rect 879 -19 883 -11
rect 742 -39 746 -35
rect 973 -1 977 3
rect 1087 -35 1091 -31
rect 900 -49 904 -45
rect 201 -69 205 -65
rect 583 -76 587 -72
rect 1160 -39 1164 -35
rect 1294 -39 1298 -35
rect 690 -69 694 -65
rect 967 -76 971 -72
rect 1388 -25 1392 -21
rect 1108 -69 1112 -65
rect 1468 -59 1472 -55
rect 1315 -73 1319 -69
rect 1536 -63 1540 -59
rect 1382 -100 1386 -96
rect 115 -110 119 -106
rect 604 -110 608 -106
rect 988 -110 992 -106
rect 1489 -93 1493 -89
rect 1403 -134 1407 -130
rect 399 -322 403 -318
rect 321 -382 325 -378
rect 32 -402 36 -398
rect 119 -410 123 -406
rect 185 -414 189 -410
rect 432 -330 436 -326
rect 456 -342 460 -338
rect 507 -358 511 -354
rect 815 -322 819 -318
rect 737 -382 741 -378
rect 848 -330 852 -326
rect 872 -342 876 -338
rect 923 -358 927 -354
rect 1265 -322 1269 -318
rect 1181 -382 1185 -378
rect 1298 -330 1302 -326
rect 1322 -342 1326 -338
rect 1373 -358 1377 -354
rect 140 -444 144 -440
rect 30 -499 34 -495
rect 321 -477 325 -473
rect 417 -459 421 -455
rect 120 -526 124 -522
rect 186 -530 190 -526
rect 450 -467 454 -463
rect 474 -479 478 -475
rect 525 -495 529 -491
rect 730 -505 734 -501
rect 833 -487 837 -483
rect 613 -547 617 -543
rect 141 -560 145 -556
rect 634 -559 638 -555
rect 679 -551 683 -547
rect 866 -495 870 -491
rect 890 -507 894 -503
rect 941 -523 945 -519
rect 1180 -474 1184 -470
rect 1283 -459 1287 -455
rect 1022 -508 1026 -504
rect 1043 -520 1047 -516
rect 1088 -512 1092 -508
rect 1316 -467 1320 -463
rect 1340 -479 1344 -475
rect 1391 -495 1395 -491
rect 1503 -500 1507 -496
rect 1532 -516 1536 -512
rect 1556 -525 1560 -521
rect 1580 -534 1584 -530
rect 1627 -508 1631 -504
rect 101 -701 105 -697
rect 122 -709 126 -705
rect 143 -717 147 -713
rect 164 -725 168 -721
rect 232 -733 236 -729
rect 371 -701 375 -697
rect 392 -710 396 -706
rect 413 -719 417 -715
rect 434 -728 438 -724
rect 502 -736 506 -732
<< metal1 >>
rect -202 147 -186 151
rect -170 147 1244 151
rect -202 122 -154 126
rect -138 122 851 126
rect -202 97 -122 101
rect -106 97 479 101
rect -202 72 -87 76
rect 47 76 216 80
rect -71 72 -61 76
rect -65 -11 -61 72
rect -14 60 59 64
rect -14 -11 -10 60
rect 55 37 59 60
rect 78 58 82 76
rect 111 58 115 76
rect 55 33 79 37
rect 88 33 92 54
rect 88 29 156 33
rect 5 25 42 29
rect 5 10 9 25
rect 38 10 42 25
rect 111 13 115 29
rect -65 -15 6 -11
rect 15 -15 19 6
rect 96 -15 100 3
rect 15 -19 100 -15
rect 38 -35 42 -19
rect 23 -107 27 -45
rect 68 -72 72 -19
rect 93 -33 134 -29
rect 152 -31 156 29
rect 179 -10 183 76
rect 212 8 216 76
rect 471 64 479 97
rect 536 76 705 80
rect 471 60 548 64
rect 212 4 309 8
rect 212 -10 216 4
rect 305 -14 309 4
rect 471 -11 479 60
rect 544 37 548 60
rect 567 58 571 76
rect 600 58 604 76
rect 544 33 568 37
rect 577 33 581 54
rect 577 29 645 33
rect 494 25 531 29
rect 494 10 498 25
rect 527 10 531 25
rect 600 13 604 29
rect 93 -51 97 -33
rect 126 -51 130 -33
rect 152 -35 180 -31
rect 189 -35 193 -14
rect 189 -39 306 -35
rect 315 -39 319 -18
rect 471 -19 495 -11
rect 504 -15 508 6
rect 585 -15 589 3
rect 504 -19 589 -15
rect 527 -35 531 -19
rect 212 -55 216 -39
rect 315 -43 351 -39
rect 315 -53 319 -43
rect 68 -76 94 -72
rect 103 -76 107 -55
rect 197 -76 201 -65
rect 103 -80 201 -76
rect 126 -96 130 -80
rect 305 -90 309 -57
rect 512 -72 516 -45
rect 192 -94 309 -90
rect 471 -80 516 -72
rect 557 -72 561 -19
rect 575 -33 623 -29
rect 641 -31 645 29
rect 668 -10 672 76
rect 701 8 705 76
rect 701 4 745 8
rect 701 -10 705 4
rect 741 -14 745 4
rect 843 -11 851 122
rect 920 76 1123 80
rect 859 60 932 64
rect 859 -11 863 60
rect 928 37 932 60
rect 951 58 955 76
rect 984 58 988 76
rect 928 33 952 37
rect 961 33 965 54
rect 961 29 1029 33
rect 878 25 915 29
rect 878 10 882 25
rect 911 10 915 25
rect 984 13 988 29
rect 582 -51 586 -33
rect 615 -51 619 -33
rect 641 -35 669 -31
rect 678 -35 682 -14
rect 678 -39 742 -35
rect 751 -39 755 -18
rect 843 -19 879 -11
rect 888 -15 892 6
rect 969 -15 973 3
rect 888 -19 973 -15
rect 911 -35 915 -19
rect 701 -55 705 -39
rect 751 -43 767 -39
rect 751 -53 755 -43
rect 557 -76 583 -72
rect 592 -76 596 -55
rect 686 -76 690 -65
rect 592 -80 690 -76
rect -202 -115 -55 -107
rect -39 -115 27 -107
rect 23 -125 27 -115
rect 111 -125 115 -106
rect 23 -129 115 -125
rect 162 -124 166 -101
rect 471 -135 479 -80
rect 512 -125 516 -80
rect 615 -96 619 -80
rect 741 -90 745 -57
rect 896 -72 900 -45
rect 681 -94 745 -90
rect 876 -80 900 -72
rect 941 -72 945 -19
rect 959 -33 1007 -29
rect 1025 -31 1029 29
rect 1086 -10 1090 76
rect 1119 8 1123 76
rect 1119 4 1163 8
rect 1119 -10 1123 4
rect 1159 -14 1163 4
rect 966 -51 970 -33
rect 999 -51 1003 -33
rect 1025 -35 1087 -31
rect 1096 -35 1100 -14
rect 1096 -39 1160 -35
rect 1169 -39 1173 -18
rect 1240 -35 1244 147
rect 1335 52 1504 56
rect 1274 36 1347 40
rect 1274 -35 1278 36
rect 1343 13 1347 36
rect 1366 34 1370 52
rect 1399 34 1403 52
rect 1343 9 1367 13
rect 1376 9 1380 30
rect 1376 5 1444 9
rect 1293 1 1330 5
rect 1293 -14 1297 1
rect 1326 -14 1330 1
rect 1399 -11 1403 5
rect 1119 -55 1123 -39
rect 1169 -43 1217 -39
rect 1240 -39 1294 -35
rect 1303 -39 1307 -18
rect 1384 -39 1388 -21
rect 1303 -43 1388 -39
rect 1169 -53 1173 -43
rect 941 -76 967 -72
rect 976 -76 980 -55
rect 1104 -76 1108 -65
rect 976 -80 1108 -76
rect 600 -125 604 -106
rect 512 -129 604 -125
rect -202 -143 273 -135
rect 289 -143 479 -135
rect 876 -163 884 -80
rect 896 -125 900 -80
rect 999 -96 1003 -80
rect 1159 -90 1163 -57
rect 1326 -59 1330 -43
rect 1099 -94 1163 -90
rect 1311 -96 1315 -69
rect 1232 -100 1315 -96
rect 1356 -96 1360 -43
rect 1381 -57 1422 -53
rect 1440 -55 1444 5
rect 1467 -34 1471 52
rect 1500 -12 1504 52
rect 1500 -16 1539 -12
rect 1500 -34 1504 -16
rect 1535 -34 1539 -16
rect 1381 -75 1385 -57
rect 1414 -75 1418 -57
rect 1440 -59 1468 -55
rect 1477 -59 1481 -38
rect 1545 -59 1549 -38
rect 1477 -63 1536 -59
rect 1545 -63 1557 -59
rect 1500 -79 1504 -63
rect 1545 -73 1549 -63
rect 1356 -100 1382 -96
rect 1391 -100 1395 -79
rect 1535 -87 1539 -77
rect 1485 -100 1489 -89
rect 1528 -91 1539 -87
rect 984 -125 988 -106
rect 896 -129 988 -125
rect -202 -171 688 -163
rect 704 -171 884 -163
rect 1232 -191 1240 -100
rect 1311 -149 1315 -100
rect 1391 -104 1489 -100
rect 1414 -120 1418 -104
rect 1399 -149 1403 -130
rect 1311 -153 1403 -149
rect -202 -194 1240 -191
rect -202 -199 1132 -194
rect 1137 -199 1240 -194
rect -101 -215 263 -207
rect -133 -232 682 -224
rect 676 -235 682 -232
rect -144 -257 1126 -249
rect 1120 -260 1126 -257
rect 184 -282 906 -278
rect 911 -282 1499 -278
rect -3 -349 95 -341
rect -3 -369 5 -349
rect -71 -377 5 -369
rect -3 -398 5 -377
rect 31 -359 67 -355
rect 31 -377 35 -359
rect 63 -362 67 -359
rect -3 -402 32 -398
rect 41 -402 45 -381
rect 59 -384 63 -363
rect 59 -388 87 -384
rect 41 -406 75 -402
rect 41 -416 45 -406
rect 31 -430 35 -420
rect 16 -434 35 -430
rect 12 -523 16 -434
rect 29 -445 52 -441
rect 29 -470 33 -445
rect 39 -495 43 -474
rect 26 -499 30 -495
rect 39 -499 51 -495
rect 39 -509 43 -499
rect 29 -523 33 -513
rect 71 -522 75 -406
rect 83 -467 87 -388
rect 91 -419 95 -349
rect 184 -363 188 -282
rect 111 -367 188 -363
rect 118 -385 122 -367
rect 151 -385 155 -367
rect 184 -385 188 -367
rect 263 -318 269 -295
rect 398 -300 402 -282
rect 453 -300 457 -282
rect 506 -300 510 -282
rect 541 -295 545 -282
rect 263 -322 399 -318
rect 263 -378 269 -322
rect 311 -339 324 -335
rect 320 -353 324 -339
rect 263 -382 321 -378
rect 330 -383 334 -357
rect 412 -354 416 -304
rect 471 -354 475 -304
rect 516 -342 520 -304
rect 516 -346 576 -342
rect 412 -358 507 -354
rect 471 -374 475 -358
rect 516 -374 520 -346
rect 115 -410 119 -406
rect 128 -410 132 -389
rect 128 -414 185 -410
rect 91 -423 108 -419
rect 104 -452 108 -423
rect 151 -430 155 -414
rect 194 -415 198 -389
rect 330 -387 385 -383
rect 330 -398 334 -387
rect 194 -419 231 -415
rect 320 -415 324 -402
rect 381 -404 385 -387
rect 398 -388 402 -378
rect 506 -388 510 -378
rect 398 -392 514 -388
rect 398 -415 402 -392
rect 541 -415 545 -378
rect 264 -419 402 -415
rect 416 -419 545 -415
rect 194 -430 198 -419
rect 136 -452 140 -440
rect 104 -456 140 -452
rect 83 -471 189 -467
rect 119 -501 123 -471
rect 152 -501 156 -471
rect 185 -501 189 -471
rect 12 -527 58 -523
rect 71 -526 120 -522
rect 129 -526 133 -505
rect 52 -567 58 -527
rect 129 -530 186 -526
rect 105 -568 109 -535
rect 152 -546 156 -530
rect 195 -531 199 -505
rect 195 -535 214 -531
rect 195 -546 199 -535
rect 137 -568 141 -556
rect 105 -572 141 -568
rect 223 -591 231 -419
rect 302 -431 324 -427
rect 298 -537 302 -431
rect 320 -445 324 -431
rect 317 -477 321 -473
rect 330 -490 334 -449
rect 320 -504 324 -494
rect 345 -504 349 -419
rect 381 -455 385 -428
rect 416 -437 420 -419
rect 471 -437 475 -419
rect 524 -437 528 -419
rect 381 -459 417 -455
rect 430 -491 434 -441
rect 489 -491 493 -441
rect 534 -479 538 -441
rect 534 -483 562 -479
rect 430 -495 525 -491
rect 320 -509 349 -504
rect 489 -511 493 -495
rect 534 -511 538 -483
rect 416 -525 420 -515
rect 524 -525 528 -515
rect 416 -529 528 -525
rect 22 -599 231 -591
rect 268 -541 302 -537
rect 268 -595 279 -541
rect 22 -721 30 -599
rect 572 -607 576 -346
rect 605 -500 609 -282
rect 676 -318 682 -295
rect 814 -300 818 -282
rect 869 -300 873 -282
rect 922 -300 926 -282
rect 676 -322 815 -318
rect 676 -378 682 -322
rect 727 -339 740 -335
rect 736 -353 740 -339
rect 676 -382 737 -378
rect 746 -383 750 -357
rect 828 -354 832 -304
rect 887 -354 891 -304
rect 932 -342 936 -304
rect 932 -346 980 -342
rect 828 -358 923 -354
rect 887 -374 891 -358
rect 932 -374 936 -346
rect 746 -387 801 -383
rect 746 -398 750 -387
rect 736 -443 740 -402
rect 797 -404 801 -387
rect 814 -388 818 -378
rect 922 -388 926 -378
rect 814 -392 926 -388
rect 814 -443 818 -392
rect 922 -419 926 -392
rect 677 -447 818 -443
rect 832 -435 907 -431
rect 718 -459 733 -455
rect 729 -473 733 -459
rect 605 -504 682 -500
rect 612 -522 616 -504
rect 645 -522 649 -504
rect 678 -522 682 -504
rect 726 -505 730 -501
rect 739 -518 743 -477
rect 588 -547 613 -543
rect 622 -547 626 -526
rect 602 -580 606 -547
rect 622 -551 679 -547
rect 614 -559 634 -555
rect 645 -567 649 -551
rect 688 -552 692 -526
rect 729 -533 733 -522
rect 761 -533 765 -447
rect 797 -483 801 -456
rect 832 -465 836 -435
rect 887 -465 891 -435
rect 912 -435 944 -431
rect 940 -465 944 -435
rect 797 -487 833 -483
rect 846 -519 850 -469
rect 905 -519 909 -469
rect 950 -507 954 -469
rect 950 -511 962 -507
rect 846 -523 941 -519
rect 729 -537 820 -533
rect 688 -556 727 -552
rect 688 -567 692 -556
rect 612 -579 616 -571
rect 678 -579 682 -571
rect 745 -579 749 -537
rect 816 -553 820 -537
rect 905 -539 909 -523
rect 950 -539 954 -511
rect 832 -553 836 -543
rect 940 -553 944 -543
rect 816 -557 944 -553
rect 612 -583 749 -579
rect 38 -615 576 -607
rect 38 -713 46 -615
rect 972 -623 980 -346
rect 1014 -461 1018 -282
rect 1120 -318 1126 -295
rect 1264 -300 1268 -282
rect 1319 -300 1323 -282
rect 1372 -283 1499 -282
rect 1372 -300 1376 -283
rect 1120 -322 1265 -318
rect 1120 -378 1126 -322
rect 1171 -339 1184 -335
rect 1180 -353 1184 -339
rect 1120 -382 1181 -378
rect 1190 -383 1194 -357
rect 1278 -354 1282 -304
rect 1337 -354 1341 -304
rect 1382 -342 1386 -304
rect 1382 -346 1430 -342
rect 1278 -358 1373 -354
rect 1337 -374 1341 -358
rect 1382 -374 1386 -346
rect 1190 -387 1251 -383
rect 1190 -398 1194 -387
rect 1180 -415 1184 -402
rect 1247 -404 1251 -387
rect 1264 -388 1268 -378
rect 1372 -388 1376 -378
rect 1264 -392 1376 -388
rect 1264 -415 1268 -392
rect 1121 -419 1268 -415
rect 1282 -419 1394 -415
rect 1014 -465 1091 -461
rect 1021 -483 1025 -465
rect 1054 -483 1058 -465
rect 1087 -483 1091 -465
rect 1006 -508 1022 -504
rect 1031 -508 1035 -487
rect 1007 -534 1011 -508
rect 1031 -512 1088 -508
rect 1023 -520 1043 -516
rect 1054 -528 1058 -512
rect 1097 -513 1101 -487
rect 1097 -517 1116 -513
rect 1097 -528 1101 -517
rect 1021 -542 1025 -532
rect 1087 -542 1091 -532
rect 1021 -546 1091 -542
rect 1112 -551 1116 -517
rect 1122 -525 1126 -419
rect 1162 -431 1183 -427
rect 1179 -445 1183 -431
rect 1176 -474 1180 -470
rect 1189 -490 1193 -449
rect 1179 -506 1183 -494
rect 1205 -506 1209 -419
rect 1247 -455 1251 -428
rect 1282 -437 1286 -419
rect 1337 -437 1341 -419
rect 1390 -437 1394 -419
rect 1247 -459 1283 -455
rect 1296 -491 1300 -441
rect 1355 -491 1359 -441
rect 1400 -479 1404 -441
rect 1400 -483 1412 -479
rect 1296 -495 1391 -491
rect 1179 -510 1209 -506
rect 1355 -511 1359 -495
rect 1400 -511 1404 -483
rect 1282 -525 1286 -515
rect 1390 -525 1394 -515
rect 1122 -529 1394 -525
rect 1122 -541 1126 -529
rect 54 -631 980 -623
rect 54 -705 62 -631
rect 1422 -639 1430 -346
rect 1495 -456 1499 -283
rect 1495 -460 1647 -456
rect 1502 -478 1506 -460
rect 1553 -478 1557 -460
rect 1594 -478 1598 -460
rect 1626 -478 1630 -460
rect 1499 -500 1503 -496
rect 1512 -504 1516 -482
rect 1573 -496 1577 -482
rect 1573 -500 1598 -496
rect 1594 -504 1598 -500
rect 1512 -508 1627 -504
rect 1499 -516 1532 -512
rect 1499 -525 1556 -521
rect 1499 -534 1580 -530
rect 1594 -540 1598 -508
rect 1636 -521 1640 -482
rect 1636 -525 1648 -521
rect 1636 -540 1640 -525
rect 1502 -552 1506 -544
rect 1626 -552 1630 -544
rect 1453 -556 1639 -552
rect 70 -647 1430 -639
rect 70 -697 78 -647
rect 100 -661 505 -657
rect 100 -679 104 -661
rect 231 -679 235 -661
rect 370 -679 374 -661
rect 501 -679 505 -661
rect 70 -701 101 -697
rect 54 -709 122 -705
rect 38 -717 143 -713
rect 22 -725 164 -721
rect 184 -729 188 -683
rect 241 -700 245 -683
rect 241 -704 253 -700
rect 361 -701 371 -697
rect 110 -733 232 -729
rect 110 -747 114 -733
rect 184 -737 188 -733
rect 157 -741 188 -737
rect 157 -747 161 -741
rect 241 -747 245 -704
rect 361 -710 392 -706
rect 361 -719 413 -715
rect 361 -728 434 -724
rect 454 -732 458 -683
rect 511 -714 515 -683
rect 511 -719 522 -714
rect 380 -736 502 -732
rect 380 -750 384 -736
rect 454 -740 458 -736
rect 427 -744 458 -740
rect 427 -750 431 -744
rect 511 -750 515 -719
rect 100 -764 104 -751
rect 133 -764 137 -751
rect 231 -764 235 -751
rect 370 -764 374 -754
rect 403 -764 407 -754
rect 501 -764 505 -754
rect 73 -768 505 -764
<< m2contact >>
rect -186 147 -170 152
rect -154 122 -138 127
rect -122 97 -106 102
rect -87 72 -71 77
rect 42 76 47 81
rect 37 29 42 34
rect 77 4 82 9
rect 4 -44 9 -39
rect 134 -33 139 -28
rect 174 10 179 15
rect 531 76 536 81
rect 526 29 531 34
rect 566 4 571 9
rect 493 -44 498 -39
rect 178 -64 183 -59
rect 187 -94 192 -89
rect 623 -33 628 -28
rect 663 10 668 15
rect 915 76 920 81
rect 910 29 915 34
rect 950 4 955 9
rect 877 -44 882 -39
rect 667 -64 672 -59
rect 92 -105 97 -100
rect 162 -101 167 -96
rect -55 -115 -39 -107
rect 162 -129 170 -124
rect 676 -94 681 -89
rect 1007 -33 1012 -28
rect 1081 10 1086 15
rect 1330 52 1335 57
rect 1325 5 1330 10
rect 1365 -20 1370 -15
rect 1085 -64 1090 -59
rect 581 -105 586 -100
rect 273 -143 289 -135
rect 1094 -94 1099 -89
rect 1292 -68 1297 -63
rect 1422 -57 1427 -52
rect 1462 -14 1467 -9
rect 1466 -88 1471 -83
rect 1528 -96 1533 -91
rect 965 -105 970 -100
rect 688 -171 704 -163
rect 1380 -129 1385 -124
rect 1132 -199 1137 -194
rect -106 -215 -101 -207
rect 263 -216 269 -207
rect -138 -232 -133 -224
rect 676 -244 682 -235
rect -149 -257 -144 -249
rect 1120 -269 1126 -260
rect 906 -282 911 -277
rect -87 -377 -71 -369
rect 63 -367 68 -362
rect 11 -434 16 -429
rect 52 -445 57 -440
rect 21 -499 26 -494
rect 51 -499 56 -494
rect 106 -367 111 -362
rect 263 -295 269 -286
rect 306 -287 311 -282
rect 540 -300 545 -295
rect 306 -339 311 -334
rect 427 -330 432 -325
rect 540 -378 545 -373
rect 108 -410 115 -405
rect 259 -419 264 -414
rect 514 -392 519 -387
rect 381 -409 386 -404
rect 117 -439 122 -434
rect 183 -439 188 -434
rect 100 -540 105 -535
rect 58 -567 63 -562
rect 214 -535 219 -530
rect 118 -555 123 -550
rect 184 -555 189 -550
rect 297 -431 302 -426
rect 312 -477 317 -472
rect 334 -484 339 -479
rect 381 -428 386 -423
rect 445 -467 450 -462
rect 562 -483 567 -478
rect 411 -529 416 -524
rect 268 -600 279 -595
rect 676 -295 682 -286
rect 722 -287 727 -282
rect 722 -339 727 -334
rect 843 -330 848 -325
rect 672 -447 677 -442
rect 797 -409 802 -404
rect 926 -419 931 -414
rect 713 -459 718 -454
rect 721 -505 726 -500
rect 743 -499 748 -494
rect 797 -456 802 -451
rect 907 -436 912 -431
rect 861 -495 866 -490
rect 962 -511 967 -506
rect 1120 -295 1126 -286
rect 1166 -287 1171 -282
rect 1355 -287 1360 -282
rect 1166 -339 1171 -334
rect 1293 -330 1298 -325
rect 1116 -419 1121 -414
rect 1247 -409 1252 -404
rect 1356 -415 1361 -410
rect 1091 -546 1096 -541
rect 1157 -431 1162 -426
rect 1171 -474 1176 -469
rect 1193 -472 1198 -467
rect 1247 -428 1252 -423
rect 1311 -467 1316 -462
rect 1412 -483 1417 -478
rect 1122 -546 1127 -541
rect 1452 -552 1457 -547
rect 268 -657 279 -652
rect 356 -701 361 -696
rect 356 -710 361 -705
rect 356 -719 361 -714
rect 356 -728 361 -723
rect 68 -768 73 -763
<< metal2 >>
rect -186 -249 -170 147
rect -154 -232 -138 122
rect -122 -215 -106 97
rect 38 85 1248 93
rect 38 81 47 85
rect -186 -257 -149 -249
rect -87 -369 -71 72
rect 38 34 42 81
rect 527 81 536 85
rect 527 34 531 81
rect 911 81 920 85
rect 911 34 915 81
rect 1244 56 1248 85
rect 1244 52 1330 56
rect 139 10 174 14
rect 628 10 663 14
rect 1012 10 1081 14
rect 1326 10 1330 52
rect 5 -53 9 -44
rect 78 -53 82 4
rect 139 -28 143 10
rect 139 -33 166 -28
rect -32 -57 82 -53
rect -55 -495 -39 -115
rect -32 -430 -28 -57
rect 78 -114 82 -57
rect 162 -96 166 -33
rect 494 -53 498 -44
rect 567 -53 571 4
rect 628 -33 632 10
rect 494 -57 571 -53
rect 878 -53 882 -44
rect 951 -53 955 4
rect 1012 -33 1016 10
rect 1427 -14 1462 -10
rect 878 -57 955 -53
rect 179 -90 183 -64
rect 179 -94 187 -90
rect 93 -114 97 -105
rect 179 -114 183 -94
rect 567 -114 571 -57
rect 668 -90 672 -64
rect 668 -94 676 -90
rect 582 -114 586 -105
rect 668 -114 672 -94
rect 951 -114 955 -57
rect 1086 -90 1090 -64
rect 1293 -77 1297 -68
rect 1366 -77 1370 -20
rect 1427 -57 1431 -14
rect 1293 -81 1370 -77
rect 1086 -94 1094 -90
rect 966 -114 970 -105
rect 1086 -114 1090 -94
rect 1366 -114 1370 -81
rect 1467 -108 1471 -88
rect 1528 -108 1532 -96
rect 78 -118 1370 -114
rect 162 -341 170 -129
rect 1366 -138 1370 -118
rect 1452 -112 1532 -108
rect 1381 -138 1385 -129
rect 1452 -138 1457 -112
rect 1366 -142 1457 -138
rect 263 -286 269 -216
rect 107 -349 170 -341
rect 107 -362 111 -349
rect 68 -367 106 -363
rect -32 -434 11 -430
rect 63 -441 69 -367
rect 57 -445 69 -441
rect 77 -410 108 -406
rect -55 -499 21 -495
rect 77 -495 81 -410
rect 118 -447 122 -439
rect 184 -447 188 -439
rect 255 -447 259 -415
rect 56 -499 81 -495
rect 92 -451 259 -447
rect 3 -536 7 -499
rect 92 -527 96 -451
rect 255 -525 259 -451
rect 273 -473 289 -143
rect 307 -334 311 -287
rect 676 -286 682 -244
rect 298 -339 306 -335
rect 371 -330 427 -326
rect 298 -426 302 -339
rect 273 -477 312 -473
rect 306 -513 310 -477
rect 371 -480 375 -330
rect 541 -373 545 -300
rect 519 -392 666 -388
rect 381 -423 385 -409
rect 658 -442 666 -392
rect 658 -447 672 -442
rect 339 -484 375 -480
rect 386 -467 445 -463
rect 386 -513 390 -467
rect 567 -483 596 -479
rect 306 -517 390 -513
rect 92 -531 114 -527
rect 255 -529 411 -525
rect 3 -540 100 -536
rect 110 -563 114 -531
rect 219 -535 247 -531
rect 119 -563 123 -555
rect 185 -563 189 -555
rect 63 -567 189 -563
rect 64 -768 68 -567
rect 239 -582 247 -535
rect 239 -587 314 -582
rect 268 -652 279 -600
rect 306 -724 314 -587
rect 592 -611 596 -483
rect 688 -501 704 -171
rect 723 -334 727 -287
rect 714 -339 722 -335
rect 787 -330 843 -326
rect 714 -454 718 -339
rect 787 -495 791 -330
rect 797 -451 801 -409
rect 907 -431 911 -282
rect 1120 -286 1126 -269
rect 931 -419 1116 -414
rect 1132 -470 1136 -199
rect 1167 -334 1171 -287
rect 1158 -339 1166 -335
rect 1237 -330 1293 -326
rect 1158 -426 1162 -339
rect 1132 -474 1171 -470
rect 1237 -468 1241 -330
rect 1247 -423 1251 -409
rect 1356 -410 1360 -287
rect 1198 -472 1241 -468
rect 1252 -467 1311 -463
rect 748 -499 791 -495
rect 802 -495 861 -491
rect 688 -505 721 -501
rect 704 -541 708 -505
rect 802 -541 806 -495
rect 967 -511 996 -507
rect 704 -545 806 -541
rect 322 -619 596 -611
rect 322 -715 330 -619
rect 988 -627 996 -511
rect 1132 -513 1136 -474
rect 1252 -513 1256 -467
rect 1417 -483 1446 -479
rect 1132 -517 1256 -513
rect 1096 -546 1122 -542
rect 336 -635 996 -627
rect 336 -706 344 -635
rect 1438 -643 1446 -483
rect 1452 -547 1457 -142
rect 348 -651 1446 -643
rect 348 -701 356 -651
rect 336 -710 356 -706
rect 322 -719 356 -715
rect 306 -728 356 -724
<< m123contact >>
rect 351 -43 359 -38
rect 767 -43 772 -38
rect 1217 -43 1225 -38
rect 1557 -64 1562 -59
rect 451 -342 456 -337
rect 469 -479 474 -474
rect 583 -547 588 -542
rect 867 -342 872 -337
rect 1317 -342 1322 -337
rect 885 -507 890 -502
rect 1001 -508 1006 -503
rect 609 -559 614 -554
rect 727 -556 732 -551
rect 601 -585 606 -580
rect 1335 -479 1340 -474
rect 1018 -520 1023 -515
rect 1007 -539 1012 -534
rect 1112 -556 1117 -551
rect 1494 -500 1499 -495
rect 1494 -516 1499 -511
rect 1494 -525 1499 -520
rect 1494 -534 1499 -529
<< metal3 >>
rect 351 -338 359 -43
rect 767 -106 771 -43
rect 676 -110 771 -106
rect 676 -157 680 -110
rect 583 -161 680 -157
rect 351 -342 451 -338
rect 351 -475 359 -342
rect 351 -479 469 -475
rect 351 -555 359 -479
rect 583 -542 587 -161
rect 1217 -179 1225 -43
rect 1557 -138 1561 -64
rect 1001 -187 1225 -179
rect 1465 -142 1561 -138
rect 767 -342 867 -338
rect 767 -503 775 -342
rect 767 -507 885 -503
rect 1001 -503 1005 -187
rect 1217 -342 1317 -338
rect 1217 -475 1225 -342
rect 1217 -479 1335 -475
rect 767 -551 775 -507
rect 351 -559 609 -555
rect 732 -556 775 -551
rect 351 -595 359 -559
rect 767 -567 775 -556
rect 999 -520 1018 -516
rect 999 -567 1003 -520
rect 767 -575 1003 -567
rect 1007 -571 1012 -539
rect 1217 -552 1225 -479
rect 1465 -496 1469 -142
rect 1465 -500 1494 -496
rect 1117 -556 1225 -552
rect 1466 -516 1494 -512
rect 1466 -571 1470 -516
rect 1007 -579 1470 -571
rect 1478 -525 1494 -521
rect 1478 -583 1482 -525
rect 606 -585 1482 -583
rect 602 -591 1482 -585
rect 1490 -595 1494 -530
rect 351 -603 1494 -595
<< labels >>
rlabel metal2 776 -498 779 -497 1 B1comp
rlabel metal2 716 -504 719 -503 1 B1
rlabel metal2 306 -476 309 -475 1 B2
rlabel metal2 361 -483 363 -482 1 B2comp
rlabel metal1 45 -498 48 -497 1 B3comp
rlabel metal1 517 -718 519 -717 1 lesser
rlabel metal1 364 -727 366 -726 1 L3
rlabel metal1 364 -718 366 -717 1 L2
rlabel metal1 364 -709 366 -708 1 L1
rlabel metal1 364 -700 366 -699 1 L0
rlabel metal1 246 -703 248 -702 1 greater
rlabel metal1 97 -700 99 -699 1 G0
rlabel metal1 97 -708 99 -707 1 G1
rlabel metal1 97 -716 99 -715 1 G2
rlabel metal1 97 -724 99 -723 1 G3
rlabel metal3 354 -571 357 -569 1 E3
rlabel metal1 339 -386 342 -385 1 A2comp
rlabel metal1 314 -381 317 -380 1 A2
rlabel metal1 321 -42 323 -41 1 E3
rlabel metal2 242 -571 244 -570 1 L3
rlabel metal1 524 -345 527 -344 1 G2
rlabel metal1 542 -482 545 -481 1 L2
rlabel metal1 729 -382 734 -380 1 A1
rlabel metal1 754 -386 759 -384 1 A1comp
rlabel metal1 940 -345 943 -344 1 G1
rlabel metal1 763 -42 765 -41 1 E2
rlabel metal1 958 -510 961 -509 1 L1
rlabel metal1 225 -571 227 -570 1 G3
rlabel metal1 -200 149 -198 151 4 A0
rlabel metal1 -200 123 -198 125 3 A1
rlabel metal2 46 87 53 91 1 VDD
rlabel metal1 -200 98 -198 100 3 A2
rlabel metal1 -201 -142 -198 -140 2 B2
rlabel metal2 -31 -56 -28 -54 1 GND
rlabel metal1 -201 -114 -199 -112 3 B3
rlabel metal1 -200 -170 -198 -168 3 B1
rlabel metal1 26 -401 29 -400 1 A3
rlabel metal1 48 -405 51 -404 1 A3comp
rlabel metal2 -2 -497 0 -496 1 B3
rlabel metal1 -201 -198 -199 -196 3 B0
rlabel metal1 -200 73 -198 75 3 A3
rlabel metal2 1163 -473 1165 -472 1 B0
rlabel metal2 1226 -472 1230 -470 1 B0comp
rlabel metal1 1552 -62 1555 -61 1 E0
rlabel metal3 1491 -537 1494 -536 1 E3
rlabel metal3 1488 -515 1491 -514 1 E1
rlabel metal3 1488 -499 1491 -498 1 E0
rlabel metal1 1643 -524 1645 -522 7 equal
rlabel metal1 1181 -42 1183 -41 1 E1
rlabel metal2 1441 -570 1444 -568 1 L0
rlabel metal1 1424 -570 1427 -568 1 G0
rlabel metal1 1174 -381 1177 -380 1 A0
rlabel metal1 1198 -386 1201 -385 1 A0comp
rlabel metal1 1390 -345 1393 -344 1 G0
rlabel metal1 1408 -482 1411 -481 1 L0
rlabel metal3 1488 -524 1491 -523 1 E2
rlabel metal1 974 -566 977 -565 1 G1
rlabel metal2 991 -565 994 -564 1 L1
rlabel metal3 763 -554 766 -553 1 E3.E2
rlabel metal3 1129 -555 1132 -554 1 E3.E2.E1
<< end >>
