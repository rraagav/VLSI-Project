magic
tech scmos
timestamp 1700498286
<< nwell >>
rect 381 98 441 122
rect 71 50 131 74
rect 308 50 368 74
rect 482 30 542 54
rect -2 2 58 26
rect 172 -18 232 6
rect 396 -11 456 13
rect 86 -59 146 -35
rect 368 -117 428 -93
rect 434 -117 462 -93
rect 527 -117 587 -93
rect 595 -117 623 -93
rect 57 -168 117 -144
rect 123 -168 151 -144
<< ntransistor >>
rect 393 61 397 69
rect 414 61 418 69
rect 83 13 87 21
rect 104 13 108 21
rect 320 13 324 21
rect 341 13 345 21
rect 10 -35 14 -27
rect 31 -35 35 -27
rect 494 -7 498 1
rect 515 -7 519 1
rect 184 -55 188 -47
rect 205 -55 209 -47
rect 408 -48 412 -40
rect 429 -48 433 -40
rect 98 -96 102 -88
rect 119 -96 123 -88
rect 380 -154 384 -146
rect 401 -154 405 -146
rect 446 -154 450 -146
rect 539 -157 543 -149
rect 560 -157 564 -149
rect 607 -157 611 -149
rect 69 -205 73 -197
rect 90 -205 94 -197
rect 135 -205 139 -197
<< ptransistor >>
rect 393 106 397 114
rect 414 106 418 114
rect 83 58 87 66
rect 104 58 108 66
rect 320 58 324 66
rect 341 58 345 66
rect 494 38 498 46
rect 515 38 519 46
rect 10 10 14 18
rect 31 10 35 18
rect 184 -10 188 -2
rect 205 -10 209 -2
rect 408 -3 412 5
rect 429 -3 433 5
rect 98 -51 102 -43
rect 119 -51 123 -43
rect 380 -109 384 -101
rect 401 -109 405 -101
rect 446 -109 450 -101
rect 539 -109 543 -101
rect 560 -109 564 -101
rect 607 -109 611 -101
rect 69 -160 73 -152
rect 90 -160 94 -152
rect 135 -160 139 -152
<< ndiffusion >>
rect 387 67 393 69
rect 387 63 388 67
rect 392 63 393 67
rect 387 61 393 63
rect 397 61 414 69
rect 418 67 435 69
rect 418 63 421 67
rect 425 63 435 67
rect 418 61 435 63
rect 77 19 83 21
rect 77 15 78 19
rect 82 15 83 19
rect 77 13 83 15
rect 87 13 104 21
rect 108 19 125 21
rect 108 15 111 19
rect 115 15 125 19
rect 108 13 125 15
rect 314 19 320 21
rect 314 15 315 19
rect 319 15 320 19
rect 314 13 320 15
rect 324 13 341 21
rect 345 19 362 21
rect 345 15 348 19
rect 352 15 362 19
rect 345 13 362 15
rect 488 -1 494 1
rect 4 -29 10 -27
rect 4 -33 5 -29
rect 9 -33 10 -29
rect 4 -35 10 -33
rect 14 -35 31 -27
rect 35 -29 52 -27
rect 35 -33 38 -29
rect 42 -33 52 -29
rect 35 -35 52 -33
rect 488 -5 489 -1
rect 493 -5 494 -1
rect 488 -7 494 -5
rect 498 -7 515 1
rect 519 -1 536 1
rect 519 -5 522 -1
rect 526 -5 536 -1
rect 519 -7 536 -5
rect 402 -42 408 -40
rect 402 -46 403 -42
rect 407 -46 408 -42
rect 178 -49 184 -47
rect 178 -53 179 -49
rect 183 -53 184 -49
rect 178 -55 184 -53
rect 188 -55 205 -47
rect 209 -49 226 -47
rect 402 -48 408 -46
rect 412 -48 429 -40
rect 433 -42 450 -40
rect 433 -46 436 -42
rect 440 -46 450 -42
rect 433 -48 450 -46
rect 209 -53 212 -49
rect 216 -53 226 -49
rect 209 -55 226 -53
rect 92 -90 98 -88
rect 92 -94 93 -90
rect 97 -94 98 -90
rect 92 -96 98 -94
rect 102 -96 119 -88
rect 123 -90 140 -88
rect 123 -94 126 -90
rect 130 -94 140 -90
rect 123 -96 140 -94
rect 374 -148 380 -146
rect 374 -152 375 -148
rect 379 -152 380 -148
rect 374 -154 380 -152
rect 384 -154 401 -146
rect 405 -148 422 -146
rect 405 -152 408 -148
rect 412 -152 422 -148
rect 405 -154 422 -152
rect 440 -148 446 -146
rect 440 -152 441 -148
rect 445 -152 446 -148
rect 440 -154 446 -152
rect 450 -148 456 -146
rect 450 -152 451 -148
rect 455 -152 456 -148
rect 450 -154 456 -152
rect 533 -151 539 -149
rect 533 -155 534 -151
rect 538 -155 539 -151
rect 533 -157 539 -155
rect 543 -151 560 -149
rect 543 -155 544 -151
rect 548 -155 560 -151
rect 543 -157 560 -155
rect 564 -151 581 -149
rect 564 -155 567 -151
rect 571 -155 581 -151
rect 564 -157 581 -155
rect 601 -151 607 -149
rect 601 -155 602 -151
rect 606 -155 607 -151
rect 601 -157 607 -155
rect 611 -151 617 -149
rect 611 -155 612 -151
rect 616 -155 617 -151
rect 611 -157 617 -155
rect 63 -199 69 -197
rect 63 -203 64 -199
rect 68 -203 69 -199
rect 63 -205 69 -203
rect 73 -205 90 -197
rect 94 -199 111 -197
rect 94 -203 97 -199
rect 101 -203 111 -199
rect 94 -205 111 -203
rect 129 -199 135 -197
rect 129 -203 130 -199
rect 134 -203 135 -199
rect 129 -205 135 -203
rect 139 -199 145 -197
rect 139 -203 140 -199
rect 144 -203 145 -199
rect 139 -205 145 -203
<< pdiffusion >>
rect 387 112 393 114
rect 387 108 388 112
rect 392 108 393 112
rect 387 106 393 108
rect 397 112 414 114
rect 397 108 398 112
rect 402 108 414 112
rect 397 106 414 108
rect 418 112 435 114
rect 418 108 421 112
rect 425 108 435 112
rect 418 106 435 108
rect 77 64 83 66
rect 77 60 78 64
rect 82 60 83 64
rect 77 58 83 60
rect 87 64 104 66
rect 87 60 88 64
rect 92 60 104 64
rect 87 58 104 60
rect 108 64 125 66
rect 108 60 111 64
rect 115 60 125 64
rect 108 58 125 60
rect 314 64 320 66
rect 314 60 315 64
rect 319 60 320 64
rect 314 58 320 60
rect 324 64 341 66
rect 324 60 325 64
rect 329 60 341 64
rect 324 58 341 60
rect 345 64 362 66
rect 345 60 348 64
rect 352 60 362 64
rect 345 58 362 60
rect 488 44 494 46
rect 488 40 489 44
rect 493 40 494 44
rect 488 38 494 40
rect 498 44 515 46
rect 498 40 499 44
rect 503 40 515 44
rect 498 38 515 40
rect 519 44 536 46
rect 519 40 522 44
rect 526 40 536 44
rect 519 38 536 40
rect 4 16 10 18
rect 4 12 5 16
rect 9 12 10 16
rect 4 10 10 12
rect 14 16 31 18
rect 14 12 15 16
rect 19 12 31 16
rect 14 10 31 12
rect 35 16 52 18
rect 35 12 38 16
rect 42 12 52 16
rect 35 10 52 12
rect 402 3 408 5
rect 402 -1 403 3
rect 407 -1 408 3
rect 178 -4 184 -2
rect 178 -8 179 -4
rect 183 -8 184 -4
rect 178 -10 184 -8
rect 188 -4 205 -2
rect 188 -8 189 -4
rect 193 -8 205 -4
rect 188 -10 205 -8
rect 209 -4 226 -2
rect 402 -3 408 -1
rect 412 3 429 5
rect 412 -1 413 3
rect 417 -1 429 3
rect 412 -3 429 -1
rect 433 3 450 5
rect 433 -1 436 3
rect 440 -1 450 3
rect 433 -3 450 -1
rect 209 -8 212 -4
rect 216 -8 226 -4
rect 209 -10 226 -8
rect 92 -45 98 -43
rect 92 -49 93 -45
rect 97 -49 98 -45
rect 92 -51 98 -49
rect 102 -45 119 -43
rect 102 -49 103 -45
rect 107 -49 119 -45
rect 102 -51 119 -49
rect 123 -45 140 -43
rect 123 -49 126 -45
rect 130 -49 140 -45
rect 123 -51 140 -49
rect 374 -103 380 -101
rect 374 -107 375 -103
rect 379 -107 380 -103
rect 374 -109 380 -107
rect 384 -103 401 -101
rect 384 -107 385 -103
rect 389 -107 401 -103
rect 384 -109 401 -107
rect 405 -103 422 -101
rect 405 -107 408 -103
rect 412 -107 422 -103
rect 405 -109 422 -107
rect 440 -103 446 -101
rect 440 -107 441 -103
rect 445 -107 446 -103
rect 440 -109 446 -107
rect 450 -103 456 -101
rect 450 -107 451 -103
rect 455 -107 456 -103
rect 450 -109 456 -107
rect 533 -103 539 -101
rect 533 -107 534 -103
rect 538 -107 539 -103
rect 533 -109 539 -107
rect 543 -109 560 -101
rect 564 -103 581 -101
rect 564 -107 569 -103
rect 573 -107 581 -103
rect 564 -109 581 -107
rect 601 -103 607 -101
rect 601 -107 602 -103
rect 606 -107 607 -103
rect 601 -109 607 -107
rect 611 -103 617 -101
rect 611 -107 612 -103
rect 616 -107 617 -103
rect 611 -109 617 -107
rect 63 -154 69 -152
rect 63 -158 64 -154
rect 68 -158 69 -154
rect 63 -160 69 -158
rect 73 -154 90 -152
rect 73 -158 74 -154
rect 78 -158 90 -154
rect 73 -160 90 -158
rect 94 -154 111 -152
rect 94 -158 97 -154
rect 101 -158 111 -154
rect 94 -160 111 -158
rect 129 -154 135 -152
rect 129 -158 130 -154
rect 134 -158 135 -154
rect 129 -160 135 -158
rect 139 -154 145 -152
rect 139 -158 140 -154
rect 144 -158 145 -154
rect 139 -160 145 -158
<< ndcontact >>
rect 388 63 392 67
rect 421 63 425 67
rect 78 15 82 19
rect 111 15 115 19
rect 315 15 319 19
rect 348 15 352 19
rect 5 -33 9 -29
rect 38 -33 42 -29
rect 489 -5 493 -1
rect 522 -5 526 -1
rect 403 -46 407 -42
rect 179 -53 183 -49
rect 436 -46 440 -42
rect 212 -53 216 -49
rect 93 -94 97 -90
rect 126 -94 130 -90
rect 375 -152 379 -148
rect 408 -152 412 -148
rect 441 -152 445 -148
rect 451 -152 455 -148
rect 534 -155 538 -151
rect 544 -155 548 -151
rect 567 -155 571 -151
rect 602 -155 606 -151
rect 612 -155 616 -151
rect 64 -203 68 -199
rect 97 -203 101 -199
rect 130 -203 134 -199
rect 140 -203 144 -199
<< pdcontact >>
rect 388 108 392 112
rect 398 108 402 112
rect 421 108 425 112
rect 78 60 82 64
rect 88 60 92 64
rect 111 60 115 64
rect 315 60 319 64
rect 325 60 329 64
rect 348 60 352 64
rect 489 40 493 44
rect 499 40 503 44
rect 522 40 526 44
rect 5 12 9 16
rect 15 12 19 16
rect 38 12 42 16
rect 403 -1 407 3
rect 179 -8 183 -4
rect 189 -8 193 -4
rect 413 -1 417 3
rect 436 -1 440 3
rect 212 -8 216 -4
rect 93 -49 97 -45
rect 103 -49 107 -45
rect 126 -49 130 -45
rect 375 -107 379 -103
rect 385 -107 389 -103
rect 408 -107 412 -103
rect 441 -107 445 -103
rect 451 -107 455 -103
rect 534 -107 538 -103
rect 569 -107 573 -103
rect 602 -107 606 -103
rect 612 -107 616 -103
rect 64 -158 68 -154
rect 74 -158 78 -154
rect 97 -158 101 -154
rect 130 -158 134 -154
rect 140 -158 144 -154
<< polysilicon >>
rect 393 114 397 117
rect 414 114 418 117
rect 393 69 397 106
rect 414 69 418 106
rect 83 66 87 69
rect 104 66 108 69
rect 320 66 324 69
rect 341 66 345 69
rect 393 58 397 61
rect 83 21 87 58
rect 104 21 108 58
rect 320 21 324 58
rect 341 21 345 58
rect 414 54 418 61
rect 494 46 498 49
rect 515 46 519 49
rect 10 18 14 21
rect 31 18 35 21
rect 83 10 87 13
rect 10 -27 14 10
rect 31 -27 35 10
rect 104 6 108 13
rect 320 10 324 13
rect 341 5 345 13
rect 408 5 412 8
rect 429 5 433 8
rect 184 -2 188 1
rect 205 -2 209 1
rect 494 1 498 38
rect 515 1 519 38
rect 10 -38 14 -35
rect 31 -43 35 -35
rect 98 -43 102 -40
rect 119 -43 123 -40
rect 184 -47 188 -10
rect 205 -47 209 -10
rect 408 -40 412 -3
rect 429 -40 433 -3
rect 494 -10 498 -7
rect 515 -15 519 -7
rect 98 -88 102 -51
rect 119 -88 123 -51
rect 408 -51 412 -48
rect 184 -58 188 -55
rect 205 -63 209 -55
rect 429 -56 433 -48
rect 98 -99 102 -96
rect 119 -104 123 -96
rect 380 -101 384 -98
rect 401 -101 405 -98
rect 446 -101 450 -98
rect 539 -101 543 -98
rect 560 -101 564 -98
rect 607 -101 611 -98
rect 380 -146 384 -109
rect 401 -146 405 -109
rect 446 -146 450 -109
rect 69 -152 73 -149
rect 90 -152 94 -149
rect 135 -152 139 -149
rect 539 -149 543 -109
rect 560 -149 564 -109
rect 607 -149 611 -109
rect 380 -157 384 -154
rect 401 -157 405 -154
rect 446 -157 450 -154
rect 539 -160 543 -157
rect 560 -160 564 -157
rect 607 -160 611 -157
rect 69 -197 73 -160
rect 90 -197 94 -160
rect 135 -197 139 -160
rect 69 -208 73 -205
rect 90 -208 94 -205
rect 135 -208 139 -205
<< polycontact >>
rect 389 87 393 91
rect 79 39 83 43
rect 316 39 320 43
rect 410 53 414 57
rect 490 19 494 23
rect 6 -9 10 -5
rect 100 5 104 9
rect 337 5 341 9
rect 180 -29 184 -25
rect 27 -43 31 -39
rect 404 -22 408 -18
rect 511 -15 515 -11
rect 94 -70 98 -66
rect 201 -63 205 -59
rect 425 -56 429 -52
rect 115 -104 119 -100
rect 376 -128 380 -124
rect 397 -140 401 -136
rect 442 -132 446 -128
rect 535 -129 539 -125
rect 556 -137 560 -133
rect 603 -145 607 -141
rect 65 -179 69 -175
rect 86 -191 90 -187
rect 131 -183 135 -179
<< metal1 >>
rect 357 130 557 134
rect 292 114 369 118
rect 47 82 247 86
rect -14 66 59 70
rect -14 -5 -10 66
rect 55 43 59 66
rect 78 64 82 82
rect 111 64 115 82
rect 55 39 79 43
rect 88 39 92 60
rect 88 35 156 39
rect 5 31 42 35
rect 5 16 9 31
rect 38 16 42 31
rect 111 19 115 35
rect -18 -9 6 -5
rect 15 -9 19 12
rect 96 -9 100 9
rect -18 -175 -14 -9
rect 15 -13 100 -9
rect 38 -29 42 -13
rect 23 -66 27 -39
rect 7 -70 27 -66
rect 68 -66 72 -13
rect 86 -27 134 -23
rect 152 -25 156 35
rect 179 -4 183 82
rect 212 -4 216 82
rect 93 -45 97 -27
rect 126 -45 130 -27
rect 152 -29 180 -25
rect 189 -31 193 -8
rect 189 -35 232 -31
rect 212 -49 216 -35
rect 68 -70 94 -66
rect 103 -70 107 -49
rect 197 -70 201 -59
rect 23 -119 27 -70
rect 103 -74 201 -70
rect 126 -90 130 -74
rect 111 -119 115 -100
rect 23 -123 115 -119
rect 27 -125 115 -123
rect 243 -132 247 82
rect 292 43 296 114
rect 365 91 369 114
rect 388 112 392 130
rect 421 112 425 130
rect 365 87 389 91
rect 398 87 402 108
rect 398 83 466 87
rect 315 79 352 83
rect 315 64 319 79
rect 348 64 352 79
rect 421 67 425 83
rect 292 39 316 43
rect 325 39 329 60
rect 406 39 410 57
rect 292 -124 296 39
rect 325 35 410 39
rect 348 19 352 35
rect 333 -18 337 9
rect 317 -22 337 -18
rect 378 -18 382 35
rect 396 21 444 25
rect 462 23 466 83
rect 489 44 493 130
rect 522 44 526 130
rect 403 3 407 21
rect 436 3 440 21
rect 462 19 490 23
rect 499 19 503 40
rect 499 15 542 19
rect 522 -1 526 15
rect 378 -22 404 -18
rect 413 -22 417 -1
rect 507 -22 511 -11
rect 333 -71 337 -22
rect 413 -26 511 -22
rect 436 -42 440 -26
rect 553 -48 557 130
rect 527 -52 557 -48
rect 421 -71 425 -52
rect 333 -75 425 -71
rect 527 -81 531 -52
rect 375 -85 606 -81
rect 375 -103 379 -85
rect 408 -103 412 -85
rect 441 -103 445 -85
rect 534 -103 538 -85
rect 602 -103 606 -85
rect 292 -128 376 -124
rect 385 -128 389 -107
rect 451 -125 455 -107
rect 385 -132 442 -128
rect 451 -129 535 -125
rect 64 -136 247 -132
rect 64 -154 68 -136
rect 97 -154 101 -136
rect 130 -154 134 -136
rect 358 -140 397 -136
rect 408 -148 412 -132
rect 451 -148 455 -129
rect 531 -137 556 -133
rect 569 -141 573 -107
rect 612 -128 616 -107
rect 612 -132 624 -128
rect 544 -145 603 -141
rect 544 -151 548 -145
rect 612 -151 616 -132
rect -18 -179 65 -175
rect 74 -179 78 -158
rect 74 -183 131 -179
rect 48 -191 86 -187
rect 97 -199 101 -183
rect 140 -184 144 -158
rect 375 -163 379 -152
rect 441 -163 445 -152
rect 368 -167 526 -163
rect 534 -167 538 -155
rect 567 -167 571 -155
rect 602 -167 606 -155
rect 522 -171 606 -167
rect 140 -188 467 -184
rect 140 -199 144 -188
rect 64 -215 68 -203
rect 130 -215 134 -203
rect 64 -219 134 -215
<< m2contact >>
rect 352 130 357 135
rect 42 82 47 87
rect 37 35 42 40
rect 77 10 82 15
rect 4 -38 9 -33
rect 134 -27 139 -22
rect 174 16 179 21
rect 232 -35 237 -30
rect 178 -58 183 -53
rect 7 -75 12 -70
rect 92 -99 97 -94
rect 347 83 352 88
rect 387 58 392 63
rect 314 10 319 15
rect 444 21 449 26
rect 484 64 489 69
rect 542 15 547 20
rect 488 -10 493 -5
rect 317 -27 322 -22
rect 402 -51 407 -46
rect 353 -141 358 -136
rect 43 -192 48 -187
rect 369 -173 374 -167
rect 467 -188 472 -183
rect 134 -219 139 -214
<< pdm12contact >>
rect 526 -137 531 -132
<< metal2 >>
rect 38 130 352 134
rect 38 40 42 130
rect 348 88 352 130
rect 449 64 484 68
rect 139 16 174 20
rect 5 -47 9 -38
rect 78 -47 82 10
rect 139 -27 143 16
rect 315 1 319 10
rect 388 1 392 58
rect 449 21 453 64
rect 547 15 563 19
rect 315 -3 392 1
rect 318 -31 322 -27
rect 237 -35 322 -31
rect -2 -51 82 -47
rect 8 -79 12 -75
rect -22 -83 12 -79
rect 8 -187 12 -83
rect 78 -108 82 -51
rect 93 -108 97 -99
rect 179 -108 183 -58
rect 78 -112 183 -108
rect 8 -191 43 -187
rect 179 -215 183 -112
rect 318 -136 322 -35
rect 388 -60 392 -3
rect 403 -60 407 -51
rect 489 -60 493 -10
rect 388 -64 493 -60
rect 318 -140 353 -136
rect 489 -169 493 -64
rect 374 -173 493 -169
rect 501 -137 526 -133
rect 403 -215 407 -173
rect 501 -183 505 -137
rect 472 -187 505 -183
rect 139 -219 407 -215
<< labels >>
rlabel metal1 292 40 294 41 1 VC
rlabel metal2 -1 -50 2 -48 1 GND
rlabel metal1 6 32 11 34 1 VDD
rlabel metal1 -18 -8 -16 -7 3 VA
rlabel metal2 -22 -82 -20 -81 3 VB
rlabel metal2 561 16 563 17 7 final_sum
rlabel metal1 616 -131 619 -129 1 final_carry
<< end >>
