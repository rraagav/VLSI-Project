* SPICE3 file created from alu.ext - technology: scmos
.include TSMC_180nm.txt

.param SUPPLY = 1
.param LAMBDA = 0.18u
.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}
.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd VDD gnd 'Supply'

Vin_S1 S1 gnd DC(0)
Vin_S0 S0 gnd DC(1)

* Vin_S0 S0 gnd PULSE(0 1 0ns 100ps 100ps 199ns 400ns)
* Vin_S1 S1 gnd PULSE(0 1 0ns 100ps 100ps 399ns 800ns)

.option scale=0.09u

M1000 VDD S0 a_200_n101# w_184_n109# CMOSP w=8 l=4
+  ad=1024 pd=480 as=136 ps=50
M1001 a_200_n146# S1 GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=480 ps=280
M1002 a_34_8# S1comp VDD w_18_0# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1003 a_34_n37# S1comp GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1004 a_34_n101# S1 VDD w_18_n109# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1005 S1comp S1 VDD w_n55_n109# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1006 a_34_8# S0comp a_34_n37# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1007 D3 a_200_n101# VDD w_250_n109# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1008 VDD S0comp a_34_8# w_18_0# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1009 a_200_8# S1comp VDD w_184_0# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1010 VDD S0comp a_34_n101# w_18_n109# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1011 a_200_n101# S1 VDD w_184_n109# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1012 D2 a_34_n101# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1013 S0comp S0 GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1014 S0comp S0 VDD w_n58_0# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1015 a_200_n101# S0 a_200_n146# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1016 D1 a_200_8# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1017 VDD S0 a_200_8# w_184_0# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1018 D1 a_200_8# VDD w_250_0# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1019 a_34_n146# S1 GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1020 D0 a_34_8# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1021 a_200_8# S0 a_200_n37# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=136 ps=50
M1022 S1comp S1 GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1023 D3 a_200_n101# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1024 D0 a_34_8# VDD w_84_0# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1025 a_200_n37# S1comp GND Gnd CMOSN w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1026 D2 a_34_n101# VDD w_84_n109# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1027 a_34_n101# S0comp a_34_n146# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
C0 S1 D0 0.09fF
C1 a_34_n101# VDD 0.03fF
C2 S0 w_184_0# 0.11fF
C3 D1 a_200_8# 0.03fF
C4 a_34_8# w_84_0# 0.11fF
C5 w_n55_n109# S1 0.11fF
C6 VDD a_34_8# 0.03fF
C7 S0comp w_n58_0# 0.03fF
C8 S1comp w_18_0# 0.11fF
C9 a_200_n101# w_250_n109# 0.11fF
C10 w_184_n109# S1 0.11fF
C11 w_84_n109# a_34_n101# 0.11fF
C12 a_200_n101# D3 0.03fF
C13 D2 S1 0.09fF
C14 w_184_0# a_200_8# 0.03fF
C15 D0 GND 0.13fF
C16 D0 w_84_0# 0.03fF
C17 w_184_0# S1comp 0.11fF
C18 VDD D0 0.08fF
C19 VDD w_n58_0# 0.03fF
C20 S1 S0comp 0.26fF
C21 w_n55_n109# VDD 0.03fF
C22 S0 w_n58_0# 0.11fF
C23 D2 GND 0.08fF
C24 w_184_n109# VDD 0.05fF
C25 S1 GND 0.35fF
C26 S1comp a_34_8# 0.03fF
C27 D2 VDD 0.03fF
C28 w_18_n109# a_34_n101# 0.03fF
C29 w_184_n109# S0 0.11fF
C30 GND S0comp 0.03fF
C31 a_34_8# w_18_0# 0.03fF
C32 D3 w_250_n109# 0.03fF
C33 S0 S1 0.19fF
C34 VDD S0comp 0.16fF
C35 D2 w_84_n109# 0.03fF
C36 a_200_n101# w_184_n109# 0.03fF
C37 a_200_n101# S1 0.03fF
C38 w_n55_n109# S1comp 0.03fF
C39 VDD GND 0.27fF
C40 S0 S0comp 0.03fF
C41 VDD w_84_0# 0.03fF
C42 S1 S1comp 0.06fF
C43 S0 GND 2.61fF
C44 w_250_0# VDD 0.03fF
C45 S0 VDD 0.25fF
C46 w_84_n109# VDD 0.03fF
C47 S1comp S0comp 0.19fF
C48 a_200_n101# VDD 0.03fF
C49 w_18_n109# S1 0.11fF
C50 GND S1comp 0.11fF
C51 VDD a_200_8# 0.03fF
C52 D0 a_34_8# 0.03fF
C53 S0comp w_18_0# 0.11fF
C54 a_200_n101# S0 0.29fF
C55 VDD S1comp 0.28fF
C56 D2 a_34_n101# 0.03fF
C57 w_18_n109# S0comp 0.11fF
C58 w_250_0# a_200_8# 0.11fF
C59 S1 a_34_n101# 0.03fF
C60 D1 GND 0.03fF
C61 S0 a_200_8# 0.29fF
C62 VDD D1 0.03fF
C63 S0 S1comp 0.19fF
C64 VDD w_18_0# 0.05fF
C65 a_34_n101# S0comp 0.29fF
C66 w_18_n109# VDD 0.05fF
C67 w_250_0# D1 0.03fF
C68 w_184_0# VDD 0.05fF
C69 D3 GND 0.03fF
C70 w_250_n109# VDD 0.03fF
C71 S0comp a_34_8# 0.29fF
C72 S1comp a_200_8# 0.03fF
C73 D3 VDD 0.03fF
C74 D3 Gnd 0.12fF
C75 D2 Gnd 0.31fF
C76 a_200_n101# Gnd 0.55fF
C77 a_34_n101# Gnd 0.55fF
C78 S1 Gnd 0.12fF
C79 GND Gnd 0.09fF
C80 D1 Gnd 0.12fF
C81 D0 Gnd 0.72fF
C82 VDD Gnd 2.80fF
C83 a_200_8# Gnd 0.55fF
C84 a_34_8# Gnd 0.55fF
C85 S0comp Gnd 0.29fF
C86 S1comp Gnd 5.74fF
C87 S0 Gnd 0.24fF
C88 w_250_n109# Gnd 0.67fF
C89 w_184_n109# Gnd 1.45fF
C90 w_84_n109# Gnd 0.67fF
C91 w_18_n109# Gnd 1.45fF
C92 w_n55_n109# Gnd 0.67fF
C93 w_250_0# Gnd 0.67fF
C94 w_184_0# Gnd 1.45fF
C95 w_84_0# Gnd 0.67fF
C96 w_18_0# Gnd 1.45fF
C97 w_n58_0# Gnd 0.67fF

.tran 1n 800n

.control
run
plot v(S0) v(S1)+2 v(D0)+4 v(D1)+6 v(D2)+8 v(D3)+10

.end
.endc