magic
tech scmos
timestamp 1700496939
<< nwell >>
rect 71 48 131 72
rect -2 0 58 24
rect 172 -20 232 4
rect 86 -61 146 -37
rect 57 -168 117 -144
rect 123 -168 151 -144
<< ntransistor >>
rect 83 11 87 19
rect 104 11 108 19
rect 10 -37 14 -29
rect 31 -37 35 -29
rect 184 -57 188 -49
rect 205 -57 209 -49
rect 98 -98 102 -90
rect 119 -98 123 -90
rect 69 -205 73 -197
rect 90 -205 94 -197
rect 135 -205 139 -197
<< ptransistor >>
rect 83 56 87 64
rect 104 56 108 64
rect 10 8 14 16
rect 31 8 35 16
rect 184 -12 188 -4
rect 205 -12 209 -4
rect 98 -53 102 -45
rect 119 -53 123 -45
rect 69 -160 73 -152
rect 90 -160 94 -152
rect 135 -160 139 -152
<< ndiffusion >>
rect 77 17 83 19
rect 77 13 78 17
rect 82 13 83 17
rect 77 11 83 13
rect 87 11 104 19
rect 108 17 125 19
rect 108 13 111 17
rect 115 13 125 17
rect 108 11 125 13
rect 4 -31 10 -29
rect 4 -35 5 -31
rect 9 -35 10 -31
rect 4 -37 10 -35
rect 14 -37 31 -29
rect 35 -31 52 -29
rect 35 -35 38 -31
rect 42 -35 52 -31
rect 35 -37 52 -35
rect 178 -51 184 -49
rect 178 -55 179 -51
rect 183 -55 184 -51
rect 178 -57 184 -55
rect 188 -57 205 -49
rect 209 -51 226 -49
rect 209 -55 212 -51
rect 216 -55 226 -51
rect 209 -57 226 -55
rect 92 -92 98 -90
rect 92 -96 93 -92
rect 97 -96 98 -92
rect 92 -98 98 -96
rect 102 -98 119 -90
rect 123 -92 140 -90
rect 123 -96 126 -92
rect 130 -96 140 -92
rect 123 -98 140 -96
rect 63 -199 69 -197
rect 63 -203 64 -199
rect 68 -203 69 -199
rect 63 -205 69 -203
rect 73 -205 90 -197
rect 94 -199 111 -197
rect 94 -203 97 -199
rect 101 -203 111 -199
rect 94 -205 111 -203
rect 129 -199 135 -197
rect 129 -203 130 -199
rect 134 -203 135 -199
rect 129 -205 135 -203
rect 139 -199 145 -197
rect 139 -203 140 -199
rect 144 -203 145 -199
rect 139 -205 145 -203
<< pdiffusion >>
rect 77 62 83 64
rect 77 58 78 62
rect 82 58 83 62
rect 77 56 83 58
rect 87 62 104 64
rect 87 58 88 62
rect 92 58 104 62
rect 87 56 104 58
rect 108 62 125 64
rect 108 58 111 62
rect 115 58 125 62
rect 108 56 125 58
rect 4 14 10 16
rect 4 10 5 14
rect 9 10 10 14
rect 4 8 10 10
rect 14 14 31 16
rect 14 10 15 14
rect 19 10 31 14
rect 14 8 31 10
rect 35 14 52 16
rect 35 10 38 14
rect 42 10 52 14
rect 35 8 52 10
rect 178 -6 184 -4
rect 178 -10 179 -6
rect 183 -10 184 -6
rect 178 -12 184 -10
rect 188 -6 205 -4
rect 188 -10 189 -6
rect 193 -10 205 -6
rect 188 -12 205 -10
rect 209 -6 226 -4
rect 209 -10 212 -6
rect 216 -10 226 -6
rect 209 -12 226 -10
rect 92 -47 98 -45
rect 92 -51 93 -47
rect 97 -51 98 -47
rect 92 -53 98 -51
rect 102 -47 119 -45
rect 102 -51 103 -47
rect 107 -51 119 -47
rect 102 -53 119 -51
rect 123 -47 140 -45
rect 123 -51 126 -47
rect 130 -51 140 -47
rect 123 -53 140 -51
rect 63 -154 69 -152
rect 63 -158 64 -154
rect 68 -158 69 -154
rect 63 -160 69 -158
rect 73 -154 90 -152
rect 73 -158 74 -154
rect 78 -158 90 -154
rect 73 -160 90 -158
rect 94 -154 111 -152
rect 94 -158 97 -154
rect 101 -158 111 -154
rect 94 -160 111 -158
rect 129 -154 135 -152
rect 129 -158 130 -154
rect 134 -158 135 -154
rect 129 -160 135 -158
rect 139 -154 145 -152
rect 139 -158 140 -154
rect 144 -158 145 -154
rect 139 -160 145 -158
<< ndcontact >>
rect 78 13 82 17
rect 111 13 115 17
rect 5 -35 9 -31
rect 38 -35 42 -31
rect 179 -55 183 -51
rect 212 -55 216 -51
rect 93 -96 97 -92
rect 126 -96 130 -92
rect 64 -203 68 -199
rect 97 -203 101 -199
rect 130 -203 134 -199
rect 140 -203 144 -199
<< pdcontact >>
rect 78 58 82 62
rect 88 58 92 62
rect 111 58 115 62
rect 5 10 9 14
rect 15 10 19 14
rect 38 10 42 14
rect 179 -10 183 -6
rect 189 -10 193 -6
rect 212 -10 216 -6
rect 93 -51 97 -47
rect 103 -51 107 -47
rect 126 -51 130 -47
rect 64 -158 68 -154
rect 74 -158 78 -154
rect 97 -158 101 -154
rect 130 -158 134 -154
rect 140 -158 144 -154
<< polysilicon >>
rect 83 64 87 67
rect 104 64 108 67
rect 83 19 87 56
rect 104 19 108 56
rect 10 16 14 19
rect 31 16 35 19
rect 83 8 87 11
rect 10 -29 14 8
rect 31 -29 35 8
rect 104 4 108 11
rect 184 -4 188 -1
rect 205 -4 209 -1
rect 10 -40 14 -37
rect 31 -45 35 -37
rect 98 -45 102 -42
rect 119 -45 123 -42
rect 184 -49 188 -12
rect 205 -49 209 -12
rect 98 -90 102 -53
rect 119 -90 123 -53
rect 184 -60 188 -57
rect 205 -65 209 -57
rect 98 -101 102 -98
rect 119 -106 123 -98
rect 69 -152 73 -149
rect 90 -152 94 -149
rect 135 -152 139 -149
rect 69 -197 73 -160
rect 90 -197 94 -160
rect 135 -197 139 -160
rect 69 -208 73 -205
rect 90 -208 94 -205
rect 135 -208 139 -205
<< polycontact >>
rect 79 37 83 41
rect 6 -11 10 -7
rect 100 3 104 7
rect 180 -31 184 -27
rect 27 -45 31 -41
rect 94 -72 98 -68
rect 201 -65 205 -61
rect 115 -106 119 -102
rect 65 -179 69 -175
rect 86 -191 90 -187
rect 131 -183 135 -179
<< metal1 >>
rect 47 80 247 84
rect -14 64 59 68
rect -14 -7 -10 64
rect 55 41 59 64
rect 78 62 82 80
rect 111 62 115 80
rect 55 37 79 41
rect 88 37 92 58
rect 88 33 156 37
rect 5 29 42 33
rect 5 14 9 29
rect 38 14 42 29
rect 111 17 115 33
rect -18 -11 6 -7
rect 15 -11 19 10
rect 96 -11 100 7
rect -18 -175 -14 -11
rect 15 -15 100 -11
rect 38 -31 42 -15
rect 23 -68 27 -41
rect 7 -72 27 -68
rect 68 -68 72 -15
rect 86 -29 134 -25
rect 152 -27 156 33
rect 179 -6 183 80
rect 212 -6 216 80
rect 93 -47 97 -29
rect 126 -47 130 -29
rect 152 -31 180 -27
rect 189 -31 193 -10
rect 189 -35 232 -31
rect 212 -51 216 -35
rect 68 -72 94 -68
rect 103 -72 107 -51
rect 197 -72 201 -61
rect 23 -121 27 -72
rect 103 -76 201 -72
rect 126 -92 130 -76
rect 111 -121 115 -102
rect 23 -125 115 -121
rect 243 -132 247 80
rect 64 -136 247 -132
rect 64 -154 68 -136
rect 97 -154 101 -136
rect 130 -154 134 -136
rect -18 -179 65 -175
rect 74 -179 78 -158
rect 74 -183 131 -179
rect 48 -191 86 -187
rect 97 -199 101 -183
rect 140 -184 144 -158
rect 140 -188 153 -184
rect 140 -199 144 -188
rect 64 -215 68 -203
rect 130 -215 134 -203
rect 64 -219 134 -215
<< m2contact >>
rect 42 80 47 85
rect 37 33 42 38
rect 77 8 82 13
rect 4 -40 9 -35
rect 134 -29 139 -24
rect 174 14 179 19
rect 232 -35 237 -30
rect 178 -60 183 -55
rect 7 -77 12 -72
rect 92 -101 97 -96
rect 43 -192 48 -187
rect 134 -219 139 -214
<< metal2 >>
rect 38 38 42 84
rect 139 14 174 18
rect 5 -49 9 -40
rect 78 -49 82 8
rect 139 -29 143 14
rect 237 -35 253 -31
rect -2 -53 82 -49
rect 8 -81 12 -77
rect -24 -85 12 -81
rect 8 -187 12 -85
rect 78 -110 82 -53
rect 93 -110 97 -101
rect 179 -110 183 -60
rect 78 -114 183 -110
rect 8 -191 43 -187
rect 179 -215 183 -114
rect 139 -219 183 -215
<< labels >>
rlabel metal2 -1 -52 2 -50 1 GND
rlabel metal1 6 30 11 32 1 VDD
rlabel metal2 250 -34 252 -33 7 half_sum
rlabel metal1 -18 -10 -16 -9 3 VA
rlabel metal2 -22 -84 -20 -83 3 VB
rlabel metal1 149 -187 151 -186 1 half_carry
<< end >>
