magic
tech scmos
timestamp 1700488856
<< nwell >>
rect 72 -6 132 18
rect 140 -6 168 18
<< ntransistor >>
rect 84 -46 88 -38
rect 105 -46 109 -38
rect 152 -46 156 -38
<< ptransistor >>
rect 84 2 88 10
rect 105 2 109 10
rect 152 2 156 10
<< ndiffusion >>
rect 78 -40 84 -38
rect 78 -44 79 -40
rect 83 -44 84 -40
rect 78 -46 84 -44
rect 88 -40 105 -38
rect 88 -44 89 -40
rect 93 -44 105 -40
rect 88 -46 105 -44
rect 109 -40 126 -38
rect 109 -44 112 -40
rect 116 -44 126 -40
rect 109 -46 126 -44
rect 146 -40 152 -38
rect 146 -44 147 -40
rect 151 -44 152 -40
rect 146 -46 152 -44
rect 156 -40 162 -38
rect 156 -44 157 -40
rect 161 -44 162 -40
rect 156 -46 162 -44
<< pdiffusion >>
rect 78 8 84 10
rect 78 4 79 8
rect 83 4 84 8
rect 78 2 84 4
rect 88 2 105 10
rect 109 8 126 10
rect 109 4 114 8
rect 118 4 126 8
rect 109 2 126 4
rect 146 8 152 10
rect 146 4 147 8
rect 151 4 152 8
rect 146 2 152 4
rect 156 8 162 10
rect 156 4 157 8
rect 161 4 162 8
rect 156 2 162 4
<< ndcontact >>
rect 79 -44 83 -40
rect 89 -44 93 -40
rect 112 -44 116 -40
rect 147 -44 151 -40
rect 157 -44 161 -40
<< pdcontact >>
rect 79 4 83 8
rect 114 4 118 8
rect 147 4 151 8
rect 157 4 161 8
<< polysilicon >>
rect 84 10 88 13
rect 105 10 109 13
rect 152 10 156 13
rect 84 -38 88 2
rect 105 -38 109 2
rect 152 -38 156 2
rect 84 -49 88 -46
rect 105 -49 109 -46
rect 152 -49 156 -46
<< polycontact >>
rect 80 -18 84 -14
rect 101 -26 105 -22
rect 148 -34 152 -30
<< metal1 >>
rect 72 26 168 30
rect 79 8 83 26
rect 147 8 151 26
rect 76 -18 80 -14
rect 76 -26 101 -22
rect 114 -30 118 4
rect 157 -17 161 4
rect 157 -21 169 -17
rect 89 -34 148 -30
rect 89 -40 93 -34
rect 157 -40 161 -21
rect 79 -56 83 -44
rect 112 -56 116 -44
rect 147 -56 151 -44
rect 72 -60 168 -56
<< labels >>
rlabel metal1 76 28 78 29 4 VDD
rlabel metal1 77 -17 79 -16 1 VA
rlabel metal1 76 -59 78 -58 2 GND
rlabel metal1 77 -25 79 -24 1 VB
rlabel metal1 161 -20 163 -19 1 Vout
<< end >>
