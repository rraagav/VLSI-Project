* SPICE3 file created from enable.ext - technology: scmos
.include TSMC_180nm.txt

.param SUPPLY = 1.8
.param LAMBDA = 0.18u
.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}
.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd VDD gnd 'Supply'

Vin_A3 A3 gnd DC(0)
Vin_A2 A2 gnd DC(1.8)
Vin_A1 A1 gnd DC(1.8)
Vin_A0 A0 gnd DC(1.8)
//7
Vin_B3 B3 gnd DC(1.8)
Vin_B2 B2 gnd DC(1.8)
Vin_B1 B1 gnd DC(1.8)
Vin_B0 B0 gnd DC(0)
//14

Vin_E E gnd DC(1.8)

.option scale=0.09u

M1000 B0out a_163_147# VDD w_213_139# CMOSP w=8 l=4
+  ad=48 pd=28 as=1856 ps=848
M1001 a_164_745# A3 GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=768 ps=448
M1002 a_161_698# E a_161_653# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=136 ps=50
M1003 a_163_194# B1 GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1004 B2out a_163_331# VDD w_213_323# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1005 a_163_331# E a_163_286# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=136 ps=50
M1006 B0out a_163_147# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1007 A3out a_164_790# VDD w_214_782# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1008 a_164_790# E a_164_745# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1009 a_161_606# A1 VDD w_145_598# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1010 a_161_561# A1 GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1011 A0out a_161_514# VDD w_211_506# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1012 B3out a_166_423# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1013 a_163_147# B0 VDD w_147_139# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1014 VDD E a_161_606# w_145_598# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1015 B2out a_163_331# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1016 a_161_606# E a_161_561# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1017 VDD E a_163_239# w_147_231# CMOSP w=8 l=4
+  ad=0 pd=0 as=136 ps=50
M1018 a_163_331# B2 VDD w_147_323# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1019 a_163_102# B0 GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1020 a_163_239# E a_163_194# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1021 A3out a_164_790# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1022 A2out a_161_698# VDD w_211_690# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1023 A0out a_161_514# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1024 a_161_514# A0 VDD w_145_506# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1025 A2out a_161_698# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1026 a_166_423# B3 VDD w_150_415# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1027 B1out a_163_239# VDD w_213_231# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1028 VDD E a_161_514# w_145_506# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1029 VDD E a_166_423# w_150_415# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1030 a_163_286# B2 GND Gnd CMOSN w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1031 B1out a_163_239# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1032 a_164_790# A3 VDD w_148_782# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1033 VDD E a_163_147# w_147_139# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1034 a_161_698# A2 VDD w_145_690# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1035 a_161_469# A0 GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1036 VDD E a_163_331# w_147_323# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1037 a_163_147# E a_163_102# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1038 a_166_378# B3 GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1039 VDD E a_164_790# w_148_782# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1040 A1out a_161_606# VDD w_211_598# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1041 a_161_653# A2 GND Gnd CMOSN w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1042 A1out a_161_606# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1043 VDD E a_161_698# w_145_690# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1044 a_161_514# E a_161_469# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1045 B3out a_166_423# VDD w_216_415# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1046 a_166_423# E a_166_378# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1047 a_163_239# B1 VDD w_147_231# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
C0 B2 E 0.19fF
C1 E A2 0.19fF
C2 a_161_514# VDD 0.03fF
C3 w_147_231# B1 0.11fF
C4 B1out w_213_231# 0.03fF
C5 A3out a_164_790# 0.03fF
C6 A0out w_211_506# 0.03fF
C7 E a_163_147# 0.29fF
C8 A2 w_145_690# 0.11fF
C9 w_145_506# E 0.11fF
C10 VDD A1 0.07fF
C11 GND B2out 0.03fF
C12 w_211_690# A2out 0.03fF
C13 a_161_514# E 0.29fF
C14 GND VDD 3.36fF
C15 A0 VDD 0.07fF
C16 w_148_782# A3 0.11fF
C17 A1out VDD 0.03fF
C18 w_150_415# a_166_423# 0.03fF
C19 B1 VDD 0.07fF
C20 E A1 0.19fF
C21 a_166_423# B3out 0.03fF
C22 w_213_323# B2out 0.03fF
C23 w_213_323# VDD 0.03fF
C24 E A0 0.19fF
C25 A3 VDD 0.07fF
C26 w_145_598# VDD 0.05fF
C27 B3out w_216_415# 0.03fF
C28 GND A2out 0.03fF
C29 E B1 0.19fF
C30 w_147_231# VDD 0.05fF
C31 a_163_147# w_147_139# 0.03fF
C32 E B0 0.19fF
C33 w_147_323# VDD 0.05fF
C34 w_148_782# VDD 0.05fF
C35 A3 a_164_790# 0.03fF
C36 E A3 0.19fF
C37 E w_145_598# 0.11fF
C38 B0out a_163_147# 0.03fF
C39 B1 a_163_239# 0.03fF
C40 a_161_514# w_211_506# 0.11fF
C41 E w_147_231# 0.11fF
C42 VDD B2out 0.03fF
C43 a_163_147# w_213_139# 0.11fF
C44 VDD a_161_698# 0.03fF
C45 E w_147_323# 0.11fF
C46 w_148_782# a_164_790# 0.03fF
C47 E w_148_782# 0.11fF
C48 w_147_231# a_163_239# 0.03fF
C49 GND B0out 0.03fF
C50 GND B3out 0.03fF
C51 E a_161_698# 0.29fF
C52 w_147_139# B0 0.11fF
C53 B2 a_163_331# 0.03fF
C54 a_164_790# VDD 0.03fF
C55 E VDD 0.43fF
C56 a_166_423# w_216_415# 0.11fF
C57 GND B1out 0.03fF
C58 a_161_698# A2out 0.03fF
C59 VDD A2out 0.03fF
C60 a_161_514# A0out 0.03fF
C61 w_211_598# a_161_606# 0.11fF
C62 w_145_690# a_161_698# 0.03fF
C63 B3 VDD 0.07fF
C64 w_145_690# VDD 0.05fF
C65 VDD a_163_239# 0.03fF
C66 E a_164_790# 0.29fF
C67 w_214_782# A3out 0.03fF
C68 GND A0out 0.03fF
C69 E B3 0.19fF
C70 E w_145_690# 0.11fF
C71 E a_163_239# 0.29fF
C72 a_161_606# A1 0.03fF
C73 w_147_139# VDD 0.05fF
C74 w_150_415# VDD 0.05fF
C75 VDD w_211_506# 0.03fF
C76 A1out a_161_606# 0.03fF
C77 B0out VDD 0.03fF
C78 B3out VDD 0.03fF
C79 w_213_323# a_163_331# 0.11fF
C80 B1out VDD 0.03fF
C81 E w_147_139# 0.11fF
C82 w_145_506# a_161_514# 0.03fF
C83 VDD w_213_139# 0.03fF
C84 w_150_415# E 0.11fF
C85 w_145_598# a_161_606# 0.03fF
C86 w_213_231# VDD 0.03fF
C87 GND A3out 0.03fF
C88 w_147_323# a_163_331# 0.03fF
C89 w_150_415# B3 0.11fF
C90 w_211_598# A1out 0.03fF
C91 w_145_506# A0 0.11fF
C92 A0out VDD 0.03fF
C93 a_161_514# A0 0.03fF
C94 a_163_331# B2out 0.03fF
C95 a_163_147# B0 0.03fF
C96 VDD a_163_331# 0.03fF
C97 B1out a_163_239# 0.03fF
C98 a_161_606# VDD 0.03fF
C99 B2 w_147_323# 0.11fF
C100 w_213_231# a_163_239# 0.11fF
C101 a_166_423# VDD 0.03fF
C102 w_216_415# VDD 0.03fF
C103 E a_163_331# 0.29fF
C104 A1out GND 0.03fF
C105 w_214_782# VDD 0.03fF
C106 E a_161_606# 0.29fF
C107 A2 a_161_698# 0.03fF
C108 w_145_598# A1 0.11fF
C109 B2 VDD 0.07fF
C110 A2 VDD 0.07fF
C111 E a_166_423# 0.29fF
C112 w_211_598# VDD 0.03fF
C113 A3out VDD 0.03fF
C114 w_211_690# a_161_698# 0.11fF
C115 w_214_782# a_164_790# 0.11fF
C116 a_163_147# VDD 0.03fF
C117 B0out w_213_139# 0.03fF
C118 w_211_690# VDD 0.03fF
C119 w_145_506# VDD 0.05fF
C120 a_166_423# B3 0.03fF
C121 B0out Gnd 0.12fF
C122 a_163_147# Gnd 0.55fF
C123 B0 Gnd 0.75fF
C124 B1out Gnd 0.12fF
C125 a_163_239# Gnd 0.55fF
C126 B1 Gnd 0.75fF
C127 B2out Gnd 0.12fF
C128 a_163_331# Gnd 0.55fF
C129 B2 Gnd 0.75fF
C130 B3out Gnd 0.11fF
C131 a_166_423# Gnd 0.55fF
C132 B3 Gnd 0.76fF
C133 A0out Gnd 0.12fF
C134 a_161_514# Gnd 0.55fF
C135 A0 Gnd 0.73fF
C136 A1out Gnd 0.12fF
C137 a_161_606# Gnd 0.55fF
C138 A1 Gnd 0.73fF
C139 A2out Gnd 0.12fF
C140 a_161_698# Gnd 0.55fF
C141 A2 Gnd 0.73fF
C142 GND Gnd 12.56fF
C143 A3out Gnd 0.12fF
C144 VDD Gnd 4.16fF
C145 a_164_790# Gnd 0.55fF
C146 E Gnd 5.80fF
C147 A3 Gnd 0.74fF
C148 w_213_139# Gnd 0.67fF
C149 w_147_139# Gnd 1.45fF
C150 w_213_231# Gnd 0.67fF
C151 w_147_231# Gnd 1.45fF
C152 w_213_323# Gnd 0.67fF
C153 w_147_323# Gnd 1.45fF
C154 w_216_415# Gnd 0.67fF
C155 w_150_415# Gnd 1.45fF
C156 w_211_506# Gnd 0.67fF
C157 w_145_506# Gnd 1.45fF
C158 w_211_598# Gnd 0.67fF
C159 w_145_598# Gnd 1.45fF
C160 w_211_690# Gnd 0.67fF
C161 w_145_690# Gnd 1.45fF
C162 w_214_782# Gnd 0.67fF
C163 w_148_782# Gnd 1.45fF

.tran 1n 800n

.control
run
plot v(A0) v(A1)+2 v(A2)+4 v(A3)+6 v(A0out)+8 v(A1out)+10 v(A2out)+12 v(A3out)+14
plot v(B0) v(B1)+2 v(B2)+4 v(B3)+6 v(B0out)+8 v(B1out)+10 v(B2out)+12 v(B3out)+14
.end
.endc