* SPICE3 file created from nand.ext - technology: scmos
.include TSMC_180nm.txt

.param SUPPLY = 1.8
.param LAMBDA = 0.18u
.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}
.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd VDD gnd 'Supply'

Vin_A VA gnd DC(1.8)
Vin_B VB gnd DC(1.8)
* Vin_VA VA gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
* Vin_VB VB gnd PULSE(0 1.8 0ns 100ps 100ps 40ns 80ns)

.option scale=0.09u

M1000 VDD VB Vout w_n2_0# CMOSP w=8 l=4
+  ad=184 pd=78 as=136 ps=50
M1001 Vout VA VDD w_n2_0# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1002 a_14_n37# VA GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=48 ps=28
M1003 Vout VB a_14_n37# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
C0 VB w_n2_0# 0.11fF
C1 VB VA 0.10fF
C2 w_n2_0# VA 0.11fF
C3 Vout VDD 0.03fF
C4 VB Vout 0.29fF
C5 Vout w_n2_0# 0.03fF
C6 VDD w_n2_0# 0.05fF
C7 Vout VA 0.03fF
C8 GND Gnd 0.07fF
C9 Vout Gnd 0.20fF
C10 VDD Gnd 0.18fF
C11 VB Gnd 0.41fF
C12 VA Gnd 0.32fF
C13 w_n2_0# Gnd 1.45fF


.tran 1n 800n

.control
run
plot v(Vout)+4 v(VB)+2 v(VA)

.end
.endc