magic
tech scmos
timestamp 1699038338
<< n_field_implant >>
rect -19 -1 19 21
<< ntransistor >>
rect -3 -32 0 -26
<< ptransistor >>
rect -3 2 0 9
<< ndiffusion >>
rect -10 -31 -9 -26
rect -4 -31 -3 -26
rect -10 -32 -3 -31
rect 0 -31 2 -26
rect 7 -31 10 -26
rect 0 -32 10 -31
<< pdiffusion >>
rect -10 4 -9 9
rect -4 4 -3 9
rect -10 2 -3 4
rect 0 4 2 9
rect 7 4 10 9
rect 0 2 10 4
<< ndcontact >>
rect -9 -31 -4 -26
rect 2 -31 7 -26
<< pdcontact >>
rect -9 4 -4 9
rect 2 4 7 9
<< polysilicon >>
rect -3 9 0 12
rect -3 -4 0 2
rect -7 -9 0 -4
rect -3 -26 0 -9
rect -3 -37 0 -32
<< polycontact >>
rect -12 -9 -7 -4
<< metal1 >>
rect -19 14 19 21
rect -9 9 -4 14
rect -18 -9 -12 -4
rect 2 -15 7 4
rect 2 -20 19 -15
rect 2 -26 7 -20
rect -9 -39 -4 -31
rect -19 -43 19 -39
<< labels >>
rlabel metal1 -16 16 -13 18 5 VDD
rlabel metal1 -17 -43 -15 -41 1 GND
<< end >>
