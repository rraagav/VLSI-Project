* SPICE3 file created from xor.ext - technology: scmos
.include TSMC_180nm.txt

.param SUPPLY = 1.8
.param LAMBDA = 0.18u
.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}
.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd VDD gnd 'Supply'

Vin_A VA gnd DC(0)
Vin_B VB gnd DC(0)

.option scale=0.09u

M1000 VDD a_14_8# a_87_56# w_71_48# CMOSP w=8 l=4
+  ad=736 pd=312 as=136 ps=50
M1001 VDD VB a_14_8# w_n2_0# CMOSP w=8 l=4
+  ad=0 pd=0 as=136 ps=50
M1002 Vout a_102_n53# a_188_n57# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=136 ps=50
M1003 a_87_56# a_14_8# a_87_11# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=136 ps=50
M1004 a_188_n57# a_87_56# GND Gnd CMOSN w=8 l=4
+  ad=0 pd=0 as=192 ps=112
M1005 a_102_n98# a_14_8# GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1006 a_102_n53# VB a_102_n98# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1007 a_87_56# VA VDD w_71_48# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1008 VDD a_102_n53# Vout w_172_n20# CMOSP w=8 l=4
+  ad=0 pd=0 as=136 ps=50
M1009 a_87_11# VA GND Gnd CMOSN w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1010 Vout a_87_56# VDD w_172_n20# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1011 a_102_n53# a_14_8# VDD w_86_n61# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1012 a_14_8# VA VDD w_n2_0# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1013 a_14_n37# VA GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1014 VDD VB a_102_n53# w_86_n61# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1015 a_14_8# VB a_14_n37# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
C0 w_n2_0# a_14_8# 0.03fF
C1 VA a_14_8# 0.03fF
C2 VDD w_86_n61# 0.05fF
C3 VDD a_14_8# 0.03fF
C4 Vout VDD 0.03fF
C5 w_71_48# a_14_8# 0.11fF
C6 a_102_n53# GND 0.09fF
C7 VB GND 0.17fF
C8 VDD w_172_n20# 0.05fF
C9 VA w_n2_0# 0.11fF
C10 a_102_n53# VB 0.10fF
C11 VDD w_n2_0# 0.05fF
C12 a_14_8# GND 0.26fF
C13 VA VDD 0.09fF
C14 w_71_48# VA 0.11fF
C15 a_102_n53# w_86_n61# 0.03fF
C16 a_87_56# a_14_8# 0.10fF
C17 Vout a_87_56# 0.03fF
C18 a_102_n53# a_14_8# 0.03fF
C19 a_102_n53# Vout 0.10fF
C20 w_86_n61# VB 0.11fF
C21 w_71_48# VDD 0.05fF
C22 a_14_8# VB 0.10fF
C23 a_87_56# w_172_n20# 0.11fF
C24 a_102_n53# w_172_n20# 0.11fF
C25 w_86_n61# a_14_8# 0.11fF
C26 w_n2_0# VB 0.11fF
C27 VA a_87_56# 0.03fF
C28 Vout w_172_n20# 0.03fF
C29 VDD a_87_56# 0.11fF
C30 w_71_48# a_87_56# 0.03fF
C31 a_102_n53# VDD 0.03fF
C32 Vout Gnd 0.21fF
C33 a_102_n53# Gnd 0.76fF
C34 GND Gnd 4.05fF
C35 VB Gnd 1.33fF
C36 a_87_56# Gnd 0.88fF
C37 VDD Gnd 0.04fF
C38 a_14_8# Gnd 1.29fF
C39 VA Gnd 1.31fF
C40 w_86_n61# Gnd 1.45fF
C41 w_172_n20# Gnd 1.45fF
C42 w_n2_0# Gnd 0.31fF
C43 w_71_48# Gnd 1.45fF

.tran 1n 800n
.control
run
plot v(VA) v(VB)+2 v(Vout)+4
.end
.endc