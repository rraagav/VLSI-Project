* SPICE3 file created from andder.ext - technology: scmos
.include TSMC_180nm.txt

.param SUPPLY = 1.8
.param LAMBDA = 0.18u
.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}
.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd VDD gnd 'Supply'

Vin_A3 A3 gnd DC(0)
Vin_A2 A2 gnd DC(1.8)
Vin_A1 A1 gnd DC(0)
Vin_A0 A0 gnd DC(1.8)

Vin_B3 B3 gnd DC(1.8)
Vin_B2 B2 gnd DC(1.8)
Vin_B1 B1 gnd DC(1.8)
Vin_B0 B0 gnd DC(1.8)

.option scale=0.09u

M1000 a_37_8# A0 VDD w_21_0# CMOSP w=8 l=4
+  ad=136 pd=50 as=928 ps=424
M1001 Ans1 a_37_n85# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=384 ps=224
M1002 a_37_n315# A3 GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1003 Ans2 a_37_n177# VDD w_87_n185# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1004 Ans0 a_37_8# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1005 a_37_n85# A1 VDD w_21_n93# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1006 a_37_n130# A1 GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1007 a_37_n270# B3 a_37_n315# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1008 VDD B0 a_37_8# w_21_0# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1009 a_37_n177# A2 VDD w_21_n185# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1010 VDD B1 a_37_n85# w_21_n93# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1011 Ans3 a_37_n270# VDD w_87_n278# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1012 a_37_n37# A0 GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1013 Ans2 a_37_n177# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1014 a_37_n85# B1 a_37_n130# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1015 VDD B2 a_37_n177# w_21_n185# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1016 a_37_8# B0 a_37_n37# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1017 a_37_n270# A3 VDD w_21_n278# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1018 a_37_n222# A2 GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1019 Ans3 a_37_n270# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1020 Ans0 a_37_8# VDD w_87_0# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1021 Ans1 a_37_n85# VDD w_87_n93# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1022 VDD B3 a_37_n270# w_21_n278# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1023 a_37_n177# B2 a_37_n222# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
C0 a_37_n85# A1 0.03fF
C1 w_21_n185# B2 0.11fF
C2 B1 A1 0.10fF
C3 VDD a_37_n270# 0.03fF
C4 A0 B0 0.10fF
C5 A0 w_21_0# 0.11fF
C6 Ans0 GND 0.03fF
C7 A0 a_37_8# 0.03fF
C8 w_87_n185# a_37_n177# 0.11fF
C9 VDD w_21_n278# 0.05fF
C10 w_21_n185# VDD 0.05fF
C11 w_21_n93# VDD 0.05fF
C12 Ans2 VDD 0.03fF
C13 VDD w_87_n93# 0.03fF
C14 a_37_n270# w_21_n278# 0.03fF
C15 B3 a_37_n270# 0.29fF
C16 a_37_n177# B2 0.29fF
C17 A2 B2 0.10fF
C18 a_37_8# w_87_0# 0.11fF
C19 Ans0 w_87_0# 0.03fF
C20 GND VDD 0.70fF
C21 A3 a_37_n270# 0.03fF
C22 B3 w_21_n278# 0.11fF
C23 a_37_n85# VDD 0.03fF
C24 VDD a_37_n177# 0.03fF
C25 A3 w_21_n278# 0.11fF
C26 A3 B3 0.10fF
C27 VDD w_87_0# 0.03fF
C28 w_21_0# B0 0.11fF
C29 Ans2 GND 0.03fF
C30 a_37_8# B0 0.29fF
C31 a_37_8# w_21_0# 0.03fF
C32 Ans0 a_37_8# 0.03fF
C33 w_87_n278# Ans3 0.03fF
C34 a_37_n85# w_21_n93# 0.03fF
C35 w_21_n185# a_37_n177# 0.03fF
C36 B1 w_21_n93# 0.11fF
C37 w_21_n185# A2 0.11fF
C38 Ans1 VDD 0.03fF
C39 Ans2 a_37_n177# 0.03fF
C40 a_37_n85# w_87_n93# 0.11fF
C41 VDD Ans3 0.03fF
C42 w_87_n185# VDD 0.03fF
C43 VDD w_21_0# 0.05fF
C44 VDD a_37_8# 0.03fF
C45 Ans0 VDD 0.03fF
C46 Ans3 a_37_n270# 0.03fF
C47 B1 a_37_n85# 0.29fF
C48 A2 a_37_n177# 0.03fF
C49 w_87_n278# VDD 0.03fF
C50 w_21_n93# A1 0.11fF
C51 Ans1 w_87_n93# 0.03fF
C52 GND Ans1 0.03fF
C53 w_87_n278# a_37_n270# 0.11fF
C54 Ans2 w_87_n185# 0.03fF
C55 GND Ans3 0.03fF
C56 a_37_n85# Ans1 0.03fF
C57 Ans3 Gnd 0.12fF
C58 a_37_n270# Gnd 0.55fF
C59 B3 Gnd 0.40fF
C60 A3 Gnd 0.19fF
C61 Ans2 Gnd 0.12fF
C62 a_37_n177# Gnd 0.55fF
C63 B2 Gnd 0.40fF
C64 A2 Gnd 0.18fF
C65 Ans1 Gnd 0.12fF
C66 a_37_n85# Gnd 0.44fF
C67 B1 Gnd 0.40fF
C68 A1 Gnd 0.25fF
C69 GND Gnd 5.25fF
C70 Ans0 Gnd 0.12fF
C71 VDD Gnd 2.54fF
C72 a_37_8# Gnd 0.44fF
C73 B0 Gnd 0.40fF
C74 A0 Gnd 0.25fF
C75 w_87_n278# Gnd 0.67fF
C76 w_21_n278# Gnd 1.45fF
C77 w_87_n185# Gnd 0.67fF
C78 w_21_n185# Gnd 1.45fF
C79 w_87_n93# Gnd 0.63fF
C80 w_21_n93# Gnd 1.45fF
C81 w_87_0# Gnd 0.63fF
C82 w_21_0# Gnd 1.45fF

.tran 1n 800n
.control
run
plot v(A0) v(A1)+2 v(A2)+4 v(A3)+6 v(B0)+8 v(B1)+10 v(B2)+12 v(B3)+14 v(Ans0)+16 v(Ans1)+18  v(Ans2)+20 v(Ans3)+22
.end
.endc