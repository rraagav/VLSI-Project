* SPICE3 file created from 4and.ext - technology: scmos
.include TSMC_180nm.txt

.param SUPPLY = 1.8
.param LAMBDA = 0.18u
.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}
.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd VDD gnd 'Supply'

Vin_VD VD gnd DC(0)
Vin_VC VC gnd DC(1.8)
Vin_VB VB gnd DC(0)
Vin_VA VA gnd DC(1.8)

.option scale=0.09u

M1000 Vout a_14_8# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=96 ps=56
M1001 Vout a_14_8# VDD w_122_0# CMOSP w=8 l=4
+  ad=48 pd=28 as=392 ps=162
M1002 a_67_n52# VC a_43_n52# Gnd CMOSN w=8 l=4
+  ad=160 pd=56 as=160 ps=56
M1003 a_14_8# VC VDD w_n2_0# CMOSP w=8 l=4
+  ad=360 pd=122 as=0 ps=0
M1004 a_14_n52# VA GND Gnd CMOSN w=8 l=4
+  ad=200 pd=66 as=0 ps=0
M1005 a_14_8# VA VDD w_n2_0# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1006 VDD VD a_14_8# w_n2_0# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1007 VDD VB a_14_8# w_n2_0# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1008 a_43_n52# VB a_14_n52# Gnd CMOSN w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1009 a_14_8# VD a_67_n52# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
C0 VC VD 0.73fF
C1 VA a_14_8# 0.03fF
C2 a_14_8# VDD 0.03fF
C3 w_n2_0# VB 0.11fF
C4 VD VA 0.10fF
C5 VC VB 0.49fF
C6 w_122_0# VDD 0.03fF
C7 VDD Vout 0.03fF
C8 Vout GND 0.03fF
C9 VD GND 0.03fF
C10 w_n2_0# VC 0.11fF
C11 VA VB 0.10fF
C12 w_n2_0# VA 0.11fF
C13 VC VA 0.10fF
C14 w_n2_0# VDD 0.08fF
C15 w_122_0# a_14_8# 0.11fF
C16 a_14_8# Vout 0.03fF
C17 VD a_14_8# 0.21fF
C18 w_122_0# Vout 0.03fF
C19 VB a_14_8# 0.35fF
C20 VD VB 0.10fF
C21 w_n2_0# a_14_8# 0.05fF
C22 VC a_14_8# 0.10fF
C23 w_n2_0# VD 0.11fF
C24 Vout Gnd 0.17fF
C25 a_14_8# Gnd 0.97fF
C26 VD Gnd 0.64fF
C27 VC Gnd 0.58fF
C28 VB Gnd 0.51fF
C29 VA Gnd 0.43fF
C30 w_122_0# Gnd 0.67fF
C31 w_n2_0# Gnd 2.80fF

.tran 1n 800n
.control
run
plot v(VA) v(VB)+2 v(VC)+4 v(VD)+6 v(Vout)+8
.end
.endc