magic
tech scmos
timestamp 1700505265
<< nwell >>
rect 71 44 131 68
rect 560 44 620 68
rect 944 44 1004 68
rect 1291 44 1351 68
rect -2 -4 58 20
rect 172 -24 232 0
rect 487 -4 547 20
rect 298 -28 326 -4
rect 661 -24 721 0
rect 871 -4 931 20
rect 734 -28 762 -4
rect 1045 -24 1105 0
rect 1218 -4 1278 20
rect 1118 -28 1146 -4
rect 1392 -24 1452 0
rect 1465 -28 1493 -4
rect 86 -65 146 -41
rect 575 -65 635 -41
rect 959 -65 1019 -41
rect 1306 -65 1366 -41
rect 391 -314 488 -290
rect 499 -314 527 -290
rect 807 -314 904 -290
rect 915 -314 943 -290
rect 1223 -314 1320 -290
rect 1331 -314 1359 -290
rect 313 -367 341 -343
rect 729 -367 757 -343
rect 1139 -367 1167 -343
rect 24 -391 52 -367
rect 111 -399 171 -375
rect 177 -399 205 -375
rect 24 -477 52 -453
rect 313 -462 341 -438
rect 409 -451 506 -427
rect 517 -451 545 -427
rect 729 -490 757 -466
rect 825 -479 922 -455
rect 933 -479 961 -455
rect 1139 -462 1167 -438
rect 1241 -451 1338 -427
rect 1349 -451 1377 -427
rect 112 -515 172 -491
rect 178 -515 206 -491
rect 1454 -509 1570 -485
rect 1576 -509 1604 -485
rect 93 -693 216 -669
rect 224 -693 252 -669
rect 363 -693 486 -669
rect 494 -693 522 -669
<< ntransistor >>
rect 83 7 87 15
rect 104 7 108 15
rect 572 7 576 15
rect 593 7 597 15
rect 10 -41 14 -33
rect 31 -41 35 -33
rect 956 7 960 15
rect 977 7 981 15
rect 499 -41 503 -33
rect 520 -41 524 -33
rect 184 -61 188 -53
rect 205 -61 209 -53
rect 310 -59 314 -51
rect 1303 7 1307 15
rect 1324 7 1328 15
rect 883 -41 887 -33
rect 904 -41 908 -33
rect 673 -61 677 -53
rect 694 -61 698 -53
rect 746 -59 750 -51
rect 1230 -41 1234 -33
rect 1251 -41 1255 -33
rect 1057 -61 1061 -53
rect 1078 -61 1082 -53
rect 1130 -59 1134 -51
rect 1404 -61 1408 -53
rect 1425 -61 1429 -53
rect 1477 -59 1481 -51
rect 98 -102 102 -94
rect 119 -102 123 -94
rect 587 -102 591 -94
rect 608 -102 612 -94
rect 971 -102 975 -94
rect 992 -102 996 -94
rect 1318 -102 1322 -94
rect 1339 -102 1343 -94
rect 36 -422 40 -414
rect 403 -380 407 -372
rect 436 -380 440 -372
rect 460 -380 464 -372
rect 511 -380 515 -372
rect 819 -380 823 -372
rect 852 -380 856 -372
rect 876 -380 880 -372
rect 927 -380 931 -372
rect 1235 -380 1239 -372
rect 1268 -380 1272 -372
rect 1292 -380 1296 -372
rect 1343 -380 1347 -372
rect 325 -404 329 -396
rect 741 -404 745 -396
rect 1151 -404 1155 -396
rect 123 -436 127 -428
rect 144 -436 148 -428
rect 189 -436 193 -428
rect 325 -499 329 -491
rect 36 -520 40 -512
rect 421 -517 425 -509
rect 454 -517 458 -509
rect 478 -517 482 -509
rect 529 -517 533 -509
rect 741 -527 745 -519
rect 1151 -499 1155 -491
rect 1253 -517 1257 -509
rect 1286 -517 1290 -509
rect 1310 -517 1314 -509
rect 1361 -517 1365 -509
rect 124 -552 128 -544
rect 145 -552 149 -544
rect 190 -552 194 -544
rect 837 -545 841 -537
rect 870 -545 874 -537
rect 894 -545 898 -537
rect 945 -545 949 -537
rect 1466 -544 1470 -536
rect 1495 -544 1499 -536
rect 1519 -544 1523 -536
rect 1543 -544 1547 -536
rect 1588 -544 1592 -536
rect 105 -753 109 -745
rect 126 -753 130 -745
rect 147 -753 151 -745
rect 168 -753 172 -745
rect 236 -753 240 -745
rect 375 -756 379 -748
rect 396 -756 400 -748
rect 417 -756 421 -748
rect 438 -756 442 -748
rect 506 -756 510 -748
<< ptransistor >>
rect 83 52 87 60
rect 104 52 108 60
rect 572 52 576 60
rect 593 52 597 60
rect 956 52 960 60
rect 977 52 981 60
rect 1303 52 1307 60
rect 1324 52 1328 60
rect 10 4 14 12
rect 31 4 35 12
rect 499 4 503 12
rect 520 4 524 12
rect 184 -16 188 -8
rect 205 -16 209 -8
rect 98 -57 102 -49
rect 119 -57 123 -49
rect 310 -20 314 -12
rect 883 4 887 12
rect 904 4 908 12
rect 673 -16 677 -8
rect 694 -16 698 -8
rect 587 -57 591 -49
rect 608 -57 612 -49
rect 746 -20 750 -12
rect 1230 4 1234 12
rect 1251 4 1255 12
rect 1057 -16 1061 -8
rect 1078 -16 1082 -8
rect 971 -57 975 -49
rect 992 -57 996 -49
rect 1130 -20 1134 -12
rect 1404 -16 1408 -8
rect 1425 -16 1429 -8
rect 1318 -57 1322 -49
rect 1339 -57 1343 -49
rect 1477 -20 1481 -12
rect 403 -306 407 -298
rect 436 -306 440 -298
rect 460 -306 464 -298
rect 511 -306 515 -298
rect 819 -306 823 -298
rect 852 -306 856 -298
rect 876 -306 880 -298
rect 927 -306 931 -298
rect 1235 -306 1239 -298
rect 1268 -306 1272 -298
rect 1292 -306 1296 -298
rect 1343 -306 1347 -298
rect 325 -359 329 -351
rect 36 -383 40 -375
rect 123 -391 127 -383
rect 144 -391 148 -383
rect 189 -391 193 -383
rect 741 -359 745 -351
rect 1151 -359 1155 -351
rect 421 -443 425 -435
rect 454 -443 458 -435
rect 478 -443 482 -435
rect 529 -443 533 -435
rect 325 -454 329 -446
rect 36 -469 40 -461
rect 124 -507 128 -499
rect 145 -507 149 -499
rect 190 -507 194 -499
rect 1253 -443 1257 -435
rect 1286 -443 1290 -435
rect 1310 -443 1314 -435
rect 1361 -443 1365 -435
rect 1151 -454 1155 -446
rect 837 -471 841 -463
rect 870 -471 874 -463
rect 894 -471 898 -463
rect 945 -471 949 -463
rect 741 -482 745 -474
rect 1466 -501 1470 -493
rect 1495 -501 1499 -493
rect 1519 -501 1523 -493
rect 1543 -501 1547 -493
rect 1588 -501 1592 -493
rect 105 -685 109 -677
rect 126 -685 130 -677
rect 147 -685 151 -677
rect 168 -685 172 -677
rect 236 -685 240 -677
rect 375 -685 379 -677
rect 396 -685 400 -677
rect 417 -685 421 -677
rect 438 -685 442 -677
rect 506 -685 510 -677
<< ndiffusion >>
rect 77 13 83 15
rect 77 9 78 13
rect 82 9 83 13
rect 77 7 83 9
rect 87 7 104 15
rect 108 13 125 15
rect 108 9 111 13
rect 115 9 125 13
rect 566 13 572 15
rect 108 7 125 9
rect 566 9 567 13
rect 571 9 572 13
rect 566 7 572 9
rect 576 7 593 15
rect 597 13 614 15
rect 597 9 600 13
rect 604 9 614 13
rect 950 13 956 15
rect 597 7 614 9
rect 4 -35 10 -33
rect 4 -39 5 -35
rect 9 -39 10 -35
rect 4 -41 10 -39
rect 14 -41 31 -33
rect 35 -35 52 -33
rect 35 -39 38 -35
rect 42 -39 52 -35
rect 35 -41 52 -39
rect 950 9 951 13
rect 955 9 956 13
rect 950 7 956 9
rect 960 7 977 15
rect 981 13 998 15
rect 981 9 984 13
rect 988 9 998 13
rect 1297 13 1303 15
rect 981 7 998 9
rect 493 -35 499 -33
rect 493 -39 494 -35
rect 498 -39 499 -35
rect 493 -41 499 -39
rect 503 -41 520 -33
rect 524 -35 541 -33
rect 524 -39 527 -35
rect 531 -39 541 -35
rect 524 -41 541 -39
rect 304 -53 310 -51
rect 178 -55 184 -53
rect 178 -59 179 -55
rect 183 -59 184 -55
rect 178 -61 184 -59
rect 188 -61 205 -53
rect 209 -55 226 -53
rect 209 -59 212 -55
rect 216 -59 226 -55
rect 304 -57 305 -53
rect 309 -57 310 -53
rect 304 -59 310 -57
rect 314 -53 320 -51
rect 314 -57 315 -53
rect 319 -57 320 -53
rect 1297 9 1298 13
rect 1302 9 1303 13
rect 1297 7 1303 9
rect 1307 7 1324 15
rect 1328 13 1345 15
rect 1328 9 1331 13
rect 1335 9 1345 13
rect 1328 7 1345 9
rect 877 -35 883 -33
rect 877 -39 878 -35
rect 882 -39 883 -35
rect 877 -41 883 -39
rect 887 -41 904 -33
rect 908 -35 925 -33
rect 908 -39 911 -35
rect 915 -39 925 -35
rect 908 -41 925 -39
rect 740 -53 746 -51
rect 667 -55 673 -53
rect 314 -59 320 -57
rect 209 -61 226 -59
rect 667 -59 668 -55
rect 672 -59 673 -55
rect 667 -61 673 -59
rect 677 -61 694 -53
rect 698 -55 715 -53
rect 698 -59 701 -55
rect 705 -59 715 -55
rect 740 -57 741 -53
rect 745 -57 746 -53
rect 740 -59 746 -57
rect 750 -53 756 -51
rect 750 -57 751 -53
rect 755 -57 756 -53
rect 1224 -35 1230 -33
rect 1224 -39 1225 -35
rect 1229 -39 1230 -35
rect 1224 -41 1230 -39
rect 1234 -41 1251 -33
rect 1255 -35 1272 -33
rect 1255 -39 1258 -35
rect 1262 -39 1272 -35
rect 1255 -41 1272 -39
rect 1124 -53 1130 -51
rect 1051 -55 1057 -53
rect 750 -59 756 -57
rect 698 -61 715 -59
rect 1051 -59 1052 -55
rect 1056 -59 1057 -55
rect 1051 -61 1057 -59
rect 1061 -61 1078 -53
rect 1082 -55 1099 -53
rect 1082 -59 1085 -55
rect 1089 -59 1099 -55
rect 1124 -57 1125 -53
rect 1129 -57 1130 -53
rect 1124 -59 1130 -57
rect 1134 -53 1140 -51
rect 1134 -57 1135 -53
rect 1139 -57 1140 -53
rect 1471 -53 1477 -51
rect 1398 -55 1404 -53
rect 1134 -59 1140 -57
rect 1082 -61 1099 -59
rect 1398 -59 1399 -55
rect 1403 -59 1404 -55
rect 1398 -61 1404 -59
rect 1408 -61 1425 -53
rect 1429 -55 1446 -53
rect 1429 -59 1432 -55
rect 1436 -59 1446 -55
rect 1471 -57 1472 -53
rect 1476 -57 1477 -53
rect 1471 -59 1477 -57
rect 1481 -53 1487 -51
rect 1481 -57 1482 -53
rect 1486 -57 1487 -53
rect 1481 -59 1487 -57
rect 1429 -61 1446 -59
rect 92 -96 98 -94
rect 92 -100 93 -96
rect 97 -100 98 -96
rect 92 -102 98 -100
rect 102 -102 119 -94
rect 123 -96 140 -94
rect 123 -100 126 -96
rect 130 -100 140 -96
rect 123 -102 140 -100
rect 581 -96 587 -94
rect 581 -100 582 -96
rect 586 -100 587 -96
rect 581 -102 587 -100
rect 591 -102 608 -94
rect 612 -96 629 -94
rect 612 -100 615 -96
rect 619 -100 629 -96
rect 612 -102 629 -100
rect 965 -96 971 -94
rect 965 -100 966 -96
rect 970 -100 971 -96
rect 965 -102 971 -100
rect 975 -102 992 -94
rect 996 -96 1013 -94
rect 996 -100 999 -96
rect 1003 -100 1013 -96
rect 996 -102 1013 -100
rect 1312 -96 1318 -94
rect 1312 -100 1313 -96
rect 1317 -100 1318 -96
rect 1312 -102 1318 -100
rect 1322 -102 1339 -94
rect 1343 -96 1360 -94
rect 1343 -100 1346 -96
rect 1350 -100 1360 -96
rect 1343 -102 1360 -100
rect -55 -115 -39 -107
rect -106 -215 -101 -207
rect -138 -232 -133 -224
rect -149 -257 -144 -249
rect 30 -416 36 -414
rect 30 -420 31 -416
rect 35 -420 36 -416
rect 30 -422 36 -420
rect 40 -416 46 -414
rect 40 -420 41 -416
rect 45 -420 46 -416
rect 40 -422 46 -420
rect 397 -374 403 -372
rect 397 -378 398 -374
rect 402 -378 403 -374
rect 397 -380 403 -378
rect 407 -380 436 -372
rect 440 -380 460 -372
rect 464 -374 482 -372
rect 464 -378 471 -374
rect 475 -378 482 -374
rect 464 -380 482 -378
rect 505 -374 511 -372
rect 505 -378 506 -374
rect 510 -378 511 -374
rect 505 -380 511 -378
rect 515 -374 521 -372
rect 515 -378 516 -374
rect 520 -378 521 -374
rect 515 -380 521 -378
rect 813 -374 819 -372
rect 813 -378 814 -374
rect 818 -378 819 -374
rect 813 -380 819 -378
rect 823 -380 852 -372
rect 856 -380 876 -372
rect 880 -374 898 -372
rect 880 -378 887 -374
rect 891 -378 898 -374
rect 880 -380 898 -378
rect 921 -374 927 -372
rect 921 -378 922 -374
rect 926 -378 927 -374
rect 921 -380 927 -378
rect 931 -374 937 -372
rect 931 -378 932 -374
rect 936 -378 937 -374
rect 931 -380 937 -378
rect 1229 -374 1235 -372
rect 1229 -378 1230 -374
rect 1234 -378 1235 -374
rect 1229 -380 1235 -378
rect 1239 -380 1268 -372
rect 1272 -380 1292 -372
rect 1296 -374 1314 -372
rect 1296 -378 1303 -374
rect 1307 -378 1314 -374
rect 1296 -380 1314 -378
rect 1337 -374 1343 -372
rect 1337 -378 1338 -374
rect 1342 -378 1343 -374
rect 1337 -380 1343 -378
rect 1347 -374 1353 -372
rect 1347 -378 1348 -374
rect 1352 -378 1353 -374
rect 1347 -380 1353 -378
rect 319 -398 325 -396
rect 319 -402 320 -398
rect 324 -402 325 -398
rect 319 -404 325 -402
rect 329 -398 335 -396
rect 329 -402 330 -398
rect 334 -402 335 -398
rect 329 -404 335 -402
rect 735 -398 741 -396
rect 735 -402 736 -398
rect 740 -402 741 -398
rect 735 -404 741 -402
rect 745 -398 751 -396
rect 745 -402 746 -398
rect 750 -402 751 -398
rect 745 -404 751 -402
rect 1145 -398 1151 -396
rect 1145 -402 1146 -398
rect 1150 -402 1151 -398
rect 1145 -404 1151 -402
rect 1155 -398 1161 -396
rect 1155 -402 1156 -398
rect 1160 -402 1161 -398
rect 1155 -404 1161 -402
rect 259 -419 264 -414
rect 1082 -419 1087 -414
rect 117 -430 123 -428
rect 117 -434 118 -430
rect 122 -434 123 -430
rect 117 -436 123 -434
rect 127 -436 144 -428
rect 148 -430 165 -428
rect 148 -434 151 -430
rect 155 -434 165 -430
rect 148 -436 165 -434
rect 183 -430 189 -428
rect 183 -434 184 -430
rect 188 -434 189 -430
rect 183 -436 189 -434
rect 193 -430 199 -428
rect 193 -434 194 -430
rect 198 -434 199 -430
rect 193 -436 199 -434
rect 319 -493 325 -491
rect 319 -497 320 -493
rect 324 -497 325 -493
rect 319 -499 325 -497
rect 329 -493 335 -491
rect 329 -497 330 -493
rect 334 -497 335 -493
rect 329 -499 335 -497
rect 30 -514 36 -512
rect 30 -518 31 -514
rect 35 -518 36 -514
rect 30 -520 36 -518
rect 40 -514 46 -512
rect 40 -518 41 -514
rect 45 -518 46 -514
rect 40 -520 46 -518
rect 100 -540 105 -535
rect 672 -447 677 -442
rect 415 -511 421 -509
rect 415 -515 416 -511
rect 420 -515 421 -511
rect 415 -517 421 -515
rect 425 -517 454 -509
rect 458 -517 478 -509
rect 482 -511 500 -509
rect 482 -515 489 -511
rect 493 -515 500 -511
rect 482 -517 500 -515
rect 523 -511 529 -509
rect 523 -515 524 -511
rect 528 -515 529 -511
rect 523 -517 529 -515
rect 533 -511 539 -509
rect 533 -515 534 -511
rect 538 -515 539 -511
rect 533 -517 539 -515
rect 735 -521 741 -519
rect 735 -525 736 -521
rect 740 -525 741 -521
rect 735 -527 741 -525
rect 745 -521 751 -519
rect 745 -525 746 -521
rect 750 -525 751 -521
rect 745 -527 751 -525
rect 1145 -493 1151 -491
rect 1145 -497 1146 -493
rect 1150 -497 1151 -493
rect 1145 -499 1151 -497
rect 1155 -493 1161 -491
rect 1155 -497 1156 -493
rect 1160 -497 1161 -493
rect 1155 -499 1161 -497
rect 1247 -511 1253 -509
rect 1247 -515 1248 -511
rect 1252 -515 1253 -511
rect 1247 -517 1253 -515
rect 1257 -517 1286 -509
rect 1290 -517 1310 -509
rect 1314 -511 1332 -509
rect 1314 -515 1321 -511
rect 1325 -515 1332 -511
rect 1314 -517 1332 -515
rect 1355 -511 1361 -509
rect 1355 -515 1356 -511
rect 1360 -515 1361 -511
rect 1355 -517 1361 -515
rect 1365 -511 1371 -509
rect 1365 -515 1366 -511
rect 1370 -515 1371 -511
rect 1365 -517 1371 -515
rect 831 -539 837 -537
rect 831 -543 832 -539
rect 836 -543 837 -539
rect 118 -546 124 -544
rect 118 -550 119 -546
rect 123 -550 124 -546
rect 118 -552 124 -550
rect 128 -552 145 -544
rect 149 -546 166 -544
rect 149 -550 152 -546
rect 156 -550 166 -546
rect 149 -552 166 -550
rect 184 -546 190 -544
rect 184 -550 185 -546
rect 189 -550 190 -546
rect 184 -552 190 -550
rect 194 -546 200 -544
rect 831 -545 837 -543
rect 841 -545 870 -537
rect 874 -545 894 -537
rect 898 -539 916 -537
rect 898 -543 905 -539
rect 909 -543 916 -539
rect 898 -545 916 -543
rect 939 -539 945 -537
rect 939 -543 940 -539
rect 944 -543 945 -539
rect 939 -545 945 -543
rect 949 -539 955 -537
rect 949 -543 950 -539
rect 954 -543 955 -539
rect 949 -545 955 -543
rect 1460 -538 1466 -536
rect 1460 -542 1461 -538
rect 1465 -542 1466 -538
rect 1460 -544 1466 -542
rect 1470 -544 1495 -536
rect 1499 -544 1519 -536
rect 1523 -544 1543 -536
rect 1547 -538 1564 -536
rect 1547 -542 1553 -538
rect 1557 -542 1564 -538
rect 1547 -544 1564 -542
rect 1582 -538 1588 -536
rect 1582 -542 1583 -538
rect 1587 -542 1588 -538
rect 1582 -544 1588 -542
rect 1592 -538 1598 -536
rect 1592 -542 1593 -538
rect 1597 -542 1598 -538
rect 1592 -544 1598 -542
rect 194 -550 195 -546
rect 199 -550 200 -546
rect 194 -552 200 -550
rect 99 -747 105 -745
rect 99 -751 100 -747
rect 104 -751 105 -747
rect 99 -753 105 -751
rect 109 -747 126 -745
rect 109 -751 110 -747
rect 114 -751 126 -747
rect 109 -753 126 -751
rect 130 -747 147 -745
rect 130 -751 133 -747
rect 137 -751 147 -747
rect 130 -753 147 -751
rect 151 -747 168 -745
rect 151 -751 157 -747
rect 161 -751 168 -747
rect 151 -753 168 -751
rect 172 -753 210 -745
rect 230 -747 236 -745
rect 230 -751 231 -747
rect 235 -751 236 -747
rect 230 -753 236 -751
rect 240 -747 246 -745
rect 240 -751 241 -747
rect 245 -751 246 -747
rect 240 -753 246 -751
rect 369 -750 375 -748
rect 369 -754 370 -750
rect 374 -754 375 -750
rect 369 -756 375 -754
rect 379 -750 396 -748
rect 379 -754 380 -750
rect 384 -754 396 -750
rect 379 -756 396 -754
rect 400 -750 417 -748
rect 400 -754 403 -750
rect 407 -754 417 -750
rect 400 -756 417 -754
rect 421 -750 438 -748
rect 421 -754 427 -750
rect 431 -754 438 -750
rect 421 -756 438 -754
rect 442 -756 480 -748
rect 500 -750 506 -748
rect 500 -754 501 -750
rect 505 -754 506 -750
rect 500 -756 506 -754
rect 510 -750 516 -748
rect 510 -754 511 -750
rect 515 -754 516 -750
rect 510 -756 516 -754
<< pdiffusion >>
rect 77 58 83 60
rect 77 54 78 58
rect 82 54 83 58
rect 77 52 83 54
rect 87 58 104 60
rect 87 54 88 58
rect 92 54 104 58
rect 87 52 104 54
rect 108 58 125 60
rect 108 54 111 58
rect 115 54 125 58
rect 108 52 125 54
rect 566 58 572 60
rect 566 54 567 58
rect 571 54 572 58
rect 566 52 572 54
rect 576 58 593 60
rect 576 54 577 58
rect 581 54 593 58
rect 576 52 593 54
rect 597 58 614 60
rect 597 54 600 58
rect 604 54 614 58
rect 597 52 614 54
rect 950 58 956 60
rect 950 54 951 58
rect 955 54 956 58
rect 950 52 956 54
rect 960 58 977 60
rect 960 54 961 58
rect 965 54 977 58
rect 960 52 977 54
rect 981 58 998 60
rect 981 54 984 58
rect 988 54 998 58
rect 981 52 998 54
rect 1297 58 1303 60
rect 1297 54 1298 58
rect 1302 54 1303 58
rect 1297 52 1303 54
rect 1307 58 1324 60
rect 1307 54 1308 58
rect 1312 54 1324 58
rect 1307 52 1324 54
rect 1328 58 1345 60
rect 1328 54 1331 58
rect 1335 54 1345 58
rect 1328 52 1345 54
rect 4 10 10 12
rect 4 6 5 10
rect 9 6 10 10
rect 4 4 10 6
rect 14 10 31 12
rect 14 6 15 10
rect 19 6 31 10
rect 14 4 31 6
rect 35 10 52 12
rect 35 6 38 10
rect 42 6 52 10
rect 493 10 499 12
rect 35 4 52 6
rect 493 6 494 10
rect 498 6 499 10
rect 493 4 499 6
rect 503 10 520 12
rect 503 6 504 10
rect 508 6 520 10
rect 503 4 520 6
rect 524 10 541 12
rect 524 6 527 10
rect 531 6 541 10
rect 877 10 883 12
rect 524 4 541 6
rect 178 -10 184 -8
rect 178 -14 179 -10
rect 183 -14 184 -10
rect 178 -16 184 -14
rect 188 -10 205 -8
rect 188 -14 189 -10
rect 193 -14 205 -10
rect 188 -16 205 -14
rect 209 -10 226 -8
rect 209 -14 212 -10
rect 216 -14 226 -10
rect 209 -16 226 -14
rect 304 -14 310 -12
rect 92 -51 98 -49
rect 92 -55 93 -51
rect 97 -55 98 -51
rect 92 -57 98 -55
rect 102 -51 119 -49
rect 102 -55 103 -51
rect 107 -55 119 -51
rect 102 -57 119 -55
rect 123 -51 140 -49
rect 123 -55 126 -51
rect 130 -55 140 -51
rect 304 -18 305 -14
rect 309 -18 310 -14
rect 304 -20 310 -18
rect 314 -14 320 -12
rect 314 -18 315 -14
rect 319 -18 320 -14
rect 314 -20 320 -18
rect 877 6 878 10
rect 882 6 883 10
rect 877 4 883 6
rect 887 10 904 12
rect 887 6 888 10
rect 892 6 904 10
rect 887 4 904 6
rect 908 10 925 12
rect 908 6 911 10
rect 915 6 925 10
rect 1224 10 1230 12
rect 908 4 925 6
rect 667 -10 673 -8
rect 667 -14 668 -10
rect 672 -14 673 -10
rect 667 -16 673 -14
rect 677 -10 694 -8
rect 677 -14 678 -10
rect 682 -14 694 -10
rect 677 -16 694 -14
rect 698 -10 715 -8
rect 698 -14 701 -10
rect 705 -14 715 -10
rect 698 -16 715 -14
rect 740 -14 746 -12
rect 581 -51 587 -49
rect 123 -57 140 -55
rect 581 -55 582 -51
rect 586 -55 587 -51
rect 581 -57 587 -55
rect 591 -51 608 -49
rect 591 -55 592 -51
rect 596 -55 608 -51
rect 591 -57 608 -55
rect 612 -51 629 -49
rect 612 -55 615 -51
rect 619 -55 629 -51
rect 740 -18 741 -14
rect 745 -18 746 -14
rect 740 -20 746 -18
rect 750 -14 756 -12
rect 750 -18 751 -14
rect 755 -18 756 -14
rect 750 -20 756 -18
rect 1224 6 1225 10
rect 1229 6 1230 10
rect 1224 4 1230 6
rect 1234 10 1251 12
rect 1234 6 1235 10
rect 1239 6 1251 10
rect 1234 4 1251 6
rect 1255 10 1272 12
rect 1255 6 1258 10
rect 1262 6 1272 10
rect 1255 4 1272 6
rect 1051 -10 1057 -8
rect 1051 -14 1052 -10
rect 1056 -14 1057 -10
rect 1051 -16 1057 -14
rect 1061 -10 1078 -8
rect 1061 -14 1062 -10
rect 1066 -14 1078 -10
rect 1061 -16 1078 -14
rect 1082 -10 1099 -8
rect 1082 -14 1085 -10
rect 1089 -14 1099 -10
rect 1082 -16 1099 -14
rect 1124 -14 1130 -12
rect 965 -51 971 -49
rect 612 -57 629 -55
rect 965 -55 966 -51
rect 970 -55 971 -51
rect 965 -57 971 -55
rect 975 -51 992 -49
rect 975 -55 976 -51
rect 980 -55 992 -51
rect 975 -57 992 -55
rect 996 -51 1013 -49
rect 996 -55 999 -51
rect 1003 -55 1013 -51
rect 1124 -18 1125 -14
rect 1129 -18 1130 -14
rect 1124 -20 1130 -18
rect 1134 -14 1140 -12
rect 1134 -18 1135 -14
rect 1139 -18 1140 -14
rect 1134 -20 1140 -18
rect 1398 -10 1404 -8
rect 1398 -14 1399 -10
rect 1403 -14 1404 -10
rect 1398 -16 1404 -14
rect 1408 -10 1425 -8
rect 1408 -14 1409 -10
rect 1413 -14 1425 -10
rect 1408 -16 1425 -14
rect 1429 -10 1446 -8
rect 1429 -14 1432 -10
rect 1436 -14 1446 -10
rect 1429 -16 1446 -14
rect 1471 -14 1477 -12
rect 1312 -51 1318 -49
rect 996 -57 1013 -55
rect 1312 -55 1313 -51
rect 1317 -55 1318 -51
rect 1312 -57 1318 -55
rect 1322 -51 1339 -49
rect 1322 -55 1323 -51
rect 1327 -55 1339 -51
rect 1322 -57 1339 -55
rect 1343 -51 1360 -49
rect 1343 -55 1346 -51
rect 1350 -55 1360 -51
rect 1471 -18 1472 -14
rect 1476 -18 1477 -14
rect 1471 -20 1477 -18
rect 1481 -14 1487 -12
rect 1481 -18 1482 -14
rect 1486 -18 1487 -14
rect 1481 -20 1487 -18
rect 1343 -57 1360 -55
rect 397 -300 403 -298
rect 397 -304 398 -300
rect 402 -304 403 -300
rect 397 -306 403 -304
rect 407 -300 436 -298
rect 407 -304 412 -300
rect 416 -304 436 -300
rect 407 -306 436 -304
rect 440 -300 460 -298
rect 440 -304 453 -300
rect 457 -304 460 -300
rect 440 -306 460 -304
rect 464 -300 482 -298
rect 464 -304 471 -300
rect 475 -304 482 -300
rect 464 -306 482 -304
rect 505 -300 511 -298
rect 505 -304 506 -300
rect 510 -304 511 -300
rect 505 -306 511 -304
rect 515 -300 521 -298
rect 515 -304 516 -300
rect 520 -304 521 -300
rect 515 -306 521 -304
rect 813 -300 819 -298
rect 813 -304 814 -300
rect 818 -304 819 -300
rect 813 -306 819 -304
rect 823 -300 852 -298
rect 823 -304 828 -300
rect 832 -304 852 -300
rect 823 -306 852 -304
rect 856 -300 876 -298
rect 856 -304 869 -300
rect 873 -304 876 -300
rect 856 -306 876 -304
rect 880 -300 898 -298
rect 880 -304 887 -300
rect 891 -304 898 -300
rect 880 -306 898 -304
rect 921 -300 927 -298
rect 921 -304 922 -300
rect 926 -304 927 -300
rect 921 -306 927 -304
rect 931 -300 937 -298
rect 931 -304 932 -300
rect 936 -304 937 -300
rect 931 -306 937 -304
rect 1229 -300 1235 -298
rect 1229 -304 1230 -300
rect 1234 -304 1235 -300
rect 1229 -306 1235 -304
rect 1239 -300 1268 -298
rect 1239 -304 1244 -300
rect 1248 -304 1268 -300
rect 1239 -306 1268 -304
rect 1272 -300 1292 -298
rect 1272 -304 1285 -300
rect 1289 -304 1292 -300
rect 1272 -306 1292 -304
rect 1296 -300 1314 -298
rect 1296 -304 1303 -300
rect 1307 -304 1314 -300
rect 1296 -306 1314 -304
rect 1337 -300 1343 -298
rect 1337 -304 1338 -300
rect 1342 -304 1343 -300
rect 1337 -306 1343 -304
rect 1347 -300 1353 -298
rect 1347 -304 1348 -300
rect 1352 -304 1353 -300
rect 1347 -306 1353 -304
rect 319 -353 325 -351
rect 319 -357 320 -353
rect 324 -357 325 -353
rect 319 -359 325 -357
rect 329 -353 335 -351
rect 329 -357 330 -353
rect 334 -357 335 -353
rect 329 -359 335 -357
rect 30 -377 36 -375
rect 30 -381 31 -377
rect 35 -381 36 -377
rect 30 -383 36 -381
rect 40 -377 46 -375
rect 40 -381 41 -377
rect 45 -381 46 -377
rect 40 -383 46 -381
rect 117 -385 123 -383
rect 117 -389 118 -385
rect 122 -389 123 -385
rect 117 -391 123 -389
rect 127 -385 144 -383
rect 127 -389 128 -385
rect 132 -389 144 -385
rect 127 -391 144 -389
rect 148 -385 165 -383
rect 148 -389 151 -385
rect 155 -389 165 -385
rect 148 -391 165 -389
rect 183 -385 189 -383
rect 183 -389 184 -385
rect 188 -389 189 -385
rect 183 -391 189 -389
rect 193 -385 199 -383
rect 193 -389 194 -385
rect 198 -389 199 -385
rect 193 -391 199 -389
rect 735 -353 741 -351
rect 735 -357 736 -353
rect 740 -357 741 -353
rect 735 -359 741 -357
rect 745 -353 751 -351
rect 745 -357 746 -353
rect 750 -357 751 -353
rect 745 -359 751 -357
rect 1145 -353 1151 -351
rect 1145 -357 1146 -353
rect 1150 -357 1151 -353
rect 1145 -359 1151 -357
rect 1155 -353 1161 -351
rect 1155 -357 1156 -353
rect 1160 -357 1161 -353
rect 1155 -359 1161 -357
rect 415 -437 421 -435
rect 415 -441 416 -437
rect 420 -441 421 -437
rect 415 -443 421 -441
rect 425 -437 454 -435
rect 425 -441 430 -437
rect 434 -441 454 -437
rect 425 -443 454 -441
rect 458 -437 478 -435
rect 458 -441 471 -437
rect 475 -441 478 -437
rect 458 -443 478 -441
rect 482 -437 500 -435
rect 482 -441 489 -437
rect 493 -441 500 -437
rect 482 -443 500 -441
rect 523 -437 529 -435
rect 523 -441 524 -437
rect 528 -441 529 -437
rect 523 -443 529 -441
rect 533 -437 539 -435
rect 533 -441 534 -437
rect 538 -441 539 -437
rect 533 -443 539 -441
rect 1247 -437 1253 -435
rect 1247 -441 1248 -437
rect 1252 -441 1253 -437
rect 319 -448 325 -446
rect 319 -452 320 -448
rect 324 -452 325 -448
rect 319 -454 325 -452
rect 329 -448 335 -446
rect 329 -452 330 -448
rect 334 -452 335 -448
rect 329 -454 335 -452
rect 30 -463 36 -461
rect 30 -467 31 -463
rect 35 -467 36 -463
rect 30 -469 36 -467
rect 40 -463 46 -461
rect 40 -467 41 -463
rect 45 -467 46 -463
rect 40 -469 46 -467
rect 118 -501 124 -499
rect 118 -505 119 -501
rect 123 -505 124 -501
rect 118 -507 124 -505
rect 128 -501 145 -499
rect 128 -505 129 -501
rect 133 -505 145 -501
rect 128 -507 145 -505
rect 149 -501 166 -499
rect 149 -505 152 -501
rect 156 -505 166 -501
rect 149 -507 166 -505
rect 184 -501 190 -499
rect 184 -505 185 -501
rect 189 -505 190 -501
rect 184 -507 190 -505
rect 194 -501 200 -499
rect 194 -505 195 -501
rect 199 -505 200 -501
rect 194 -507 200 -505
rect 1247 -443 1253 -441
rect 1257 -437 1286 -435
rect 1257 -441 1262 -437
rect 1266 -441 1286 -437
rect 1257 -443 1286 -441
rect 1290 -437 1310 -435
rect 1290 -441 1303 -437
rect 1307 -441 1310 -437
rect 1290 -443 1310 -441
rect 1314 -437 1332 -435
rect 1314 -441 1321 -437
rect 1325 -441 1332 -437
rect 1314 -443 1332 -441
rect 1355 -437 1361 -435
rect 1355 -441 1356 -437
rect 1360 -441 1361 -437
rect 1355 -443 1361 -441
rect 1365 -437 1371 -435
rect 1365 -441 1366 -437
rect 1370 -441 1371 -437
rect 1365 -443 1371 -441
rect 1145 -448 1151 -446
rect 1145 -452 1146 -448
rect 1150 -452 1151 -448
rect 1145 -454 1151 -452
rect 1155 -448 1161 -446
rect 1155 -452 1156 -448
rect 1160 -452 1161 -448
rect 1155 -454 1161 -452
rect 831 -465 837 -463
rect 831 -469 832 -465
rect 836 -469 837 -465
rect 831 -471 837 -469
rect 841 -465 870 -463
rect 841 -469 846 -465
rect 850 -469 870 -465
rect 841 -471 870 -469
rect 874 -465 894 -463
rect 874 -469 887 -465
rect 891 -469 894 -465
rect 874 -471 894 -469
rect 898 -465 916 -463
rect 898 -469 905 -465
rect 909 -469 916 -465
rect 898 -471 916 -469
rect 939 -465 945 -463
rect 939 -469 940 -465
rect 944 -469 945 -465
rect 939 -471 945 -469
rect 949 -465 955 -463
rect 949 -469 950 -465
rect 954 -469 955 -465
rect 949 -471 955 -469
rect 735 -476 741 -474
rect 735 -480 736 -476
rect 740 -480 741 -476
rect 735 -482 741 -480
rect 745 -476 751 -474
rect 745 -480 746 -476
rect 750 -480 751 -476
rect 745 -482 751 -480
rect 1460 -495 1466 -493
rect 1460 -499 1461 -495
rect 1465 -499 1466 -495
rect 1460 -501 1466 -499
rect 1470 -495 1495 -493
rect 1470 -499 1471 -495
rect 1475 -499 1495 -495
rect 1470 -501 1495 -499
rect 1499 -495 1519 -493
rect 1499 -499 1512 -495
rect 1516 -499 1519 -495
rect 1499 -501 1519 -499
rect 1523 -495 1543 -493
rect 1523 -499 1532 -495
rect 1536 -499 1543 -495
rect 1523 -501 1543 -499
rect 1547 -495 1564 -493
rect 1547 -499 1553 -495
rect 1557 -499 1564 -495
rect 1547 -501 1564 -499
rect 1582 -495 1588 -493
rect 1582 -499 1583 -495
rect 1587 -499 1588 -495
rect 1582 -501 1588 -499
rect 1592 -495 1598 -493
rect 1592 -499 1593 -495
rect 1597 -499 1598 -495
rect 1592 -501 1598 -499
rect 99 -679 105 -677
rect 99 -683 100 -679
rect 104 -683 105 -679
rect 99 -685 105 -683
rect 109 -685 126 -677
rect 130 -685 147 -677
rect 151 -685 168 -677
rect 172 -679 210 -677
rect 172 -683 184 -679
rect 188 -683 210 -679
rect 172 -685 210 -683
rect 230 -679 236 -677
rect 230 -683 231 -679
rect 235 -683 236 -679
rect 230 -685 236 -683
rect 240 -679 246 -677
rect 240 -683 241 -679
rect 245 -683 246 -679
rect 240 -685 246 -683
rect 369 -679 375 -677
rect 369 -683 370 -679
rect 374 -683 375 -679
rect 369 -685 375 -683
rect 379 -685 396 -677
rect 400 -685 417 -677
rect 421 -685 438 -677
rect 442 -679 480 -677
rect 442 -683 454 -679
rect 458 -683 480 -679
rect 442 -685 480 -683
rect 500 -679 506 -677
rect 500 -683 501 -679
rect 505 -683 506 -679
rect 500 -685 506 -683
rect 510 -679 516 -677
rect 510 -683 511 -679
rect 515 -683 516 -679
rect 510 -685 516 -683
<< ndcontact >>
rect 78 9 82 13
rect 111 9 115 13
rect 567 9 571 13
rect 600 9 604 13
rect 5 -39 9 -35
rect 38 -39 42 -35
rect 951 9 955 13
rect 984 9 988 13
rect 494 -39 498 -35
rect 527 -39 531 -35
rect 179 -59 183 -55
rect 212 -59 216 -55
rect 305 -57 309 -53
rect 315 -57 319 -53
rect 1298 9 1302 13
rect 1331 9 1335 13
rect 878 -39 882 -35
rect 911 -39 915 -35
rect 668 -59 672 -55
rect 701 -59 705 -55
rect 741 -57 745 -53
rect 751 -57 755 -53
rect 1225 -39 1229 -35
rect 1258 -39 1262 -35
rect 1052 -59 1056 -55
rect 1085 -59 1089 -55
rect 1125 -57 1129 -53
rect 1135 -57 1139 -53
rect 1399 -59 1403 -55
rect 1432 -59 1436 -55
rect 1472 -57 1476 -53
rect 1482 -57 1486 -53
rect 93 -100 97 -96
rect 126 -100 130 -96
rect 582 -100 586 -96
rect 615 -100 619 -96
rect 966 -100 970 -96
rect 999 -100 1003 -96
rect 1313 -100 1317 -96
rect 1346 -100 1350 -96
rect 31 -420 35 -416
rect 41 -420 45 -416
rect 398 -378 402 -374
rect 471 -378 475 -374
rect 506 -378 510 -374
rect 516 -378 520 -374
rect 814 -378 818 -374
rect 887 -378 891 -374
rect 922 -378 926 -374
rect 932 -378 936 -374
rect 1230 -378 1234 -374
rect 1303 -378 1307 -374
rect 1338 -378 1342 -374
rect 1348 -378 1352 -374
rect 320 -402 324 -398
rect 330 -402 334 -398
rect 736 -402 740 -398
rect 746 -402 750 -398
rect 1146 -402 1150 -398
rect 1156 -402 1160 -398
rect 118 -434 122 -430
rect 151 -434 155 -430
rect 184 -434 188 -430
rect 194 -434 198 -430
rect 320 -497 324 -493
rect 330 -497 334 -493
rect 31 -518 35 -514
rect 41 -518 45 -514
rect 416 -515 420 -511
rect 489 -515 493 -511
rect 524 -515 528 -511
rect 534 -515 538 -511
rect 736 -525 740 -521
rect 746 -525 750 -521
rect 1146 -497 1150 -493
rect 1156 -497 1160 -493
rect 1248 -515 1252 -511
rect 1321 -515 1325 -511
rect 1356 -515 1360 -511
rect 1366 -515 1370 -511
rect 832 -543 836 -539
rect 119 -550 123 -546
rect 152 -550 156 -546
rect 185 -550 189 -546
rect 905 -543 909 -539
rect 940 -543 944 -539
rect 950 -543 954 -539
rect 1461 -542 1465 -538
rect 1553 -542 1557 -538
rect 1583 -542 1587 -538
rect 1593 -542 1597 -538
rect 195 -550 199 -546
rect 100 -751 104 -747
rect 110 -751 114 -747
rect 133 -751 137 -747
rect 157 -751 161 -747
rect 231 -751 235 -747
rect 241 -751 245 -747
rect 370 -754 374 -750
rect 380 -754 384 -750
rect 403 -754 407 -750
rect 427 -754 431 -750
rect 501 -754 505 -750
rect 511 -754 515 -750
<< pdcontact >>
rect 78 54 82 58
rect 88 54 92 58
rect 111 54 115 58
rect 567 54 571 58
rect 577 54 581 58
rect 600 54 604 58
rect 951 54 955 58
rect 961 54 965 58
rect 984 54 988 58
rect 1298 54 1302 58
rect 1308 54 1312 58
rect 1331 54 1335 58
rect 5 6 9 10
rect 15 6 19 10
rect 38 6 42 10
rect 494 6 498 10
rect 504 6 508 10
rect 527 6 531 10
rect 179 -14 183 -10
rect 189 -14 193 -10
rect 212 -14 216 -10
rect 93 -55 97 -51
rect 103 -55 107 -51
rect 126 -55 130 -51
rect 305 -18 309 -14
rect 315 -18 319 -14
rect 878 6 882 10
rect 888 6 892 10
rect 911 6 915 10
rect 668 -14 672 -10
rect 678 -14 682 -10
rect 701 -14 705 -10
rect 582 -55 586 -51
rect 592 -55 596 -51
rect 615 -55 619 -51
rect 741 -18 745 -14
rect 751 -18 755 -14
rect 1225 6 1229 10
rect 1235 6 1239 10
rect 1258 6 1262 10
rect 1052 -14 1056 -10
rect 1062 -14 1066 -10
rect 1085 -14 1089 -10
rect 966 -55 970 -51
rect 976 -55 980 -51
rect 999 -55 1003 -51
rect 1125 -18 1129 -14
rect 1135 -18 1139 -14
rect 1399 -14 1403 -10
rect 1409 -14 1413 -10
rect 1432 -14 1436 -10
rect 1313 -55 1317 -51
rect 1323 -55 1327 -51
rect 1346 -55 1350 -51
rect 1472 -18 1476 -14
rect 1482 -18 1486 -14
rect 398 -304 402 -300
rect 412 -304 416 -300
rect 453 -304 457 -300
rect 471 -304 475 -300
rect 506 -304 510 -300
rect 516 -304 520 -300
rect 814 -304 818 -300
rect 828 -304 832 -300
rect 869 -304 873 -300
rect 887 -304 891 -300
rect 922 -304 926 -300
rect 932 -304 936 -300
rect 1230 -304 1234 -300
rect 1244 -304 1248 -300
rect 1285 -304 1289 -300
rect 1303 -304 1307 -300
rect 1338 -304 1342 -300
rect 1348 -304 1352 -300
rect 320 -357 324 -353
rect 330 -357 334 -353
rect 31 -381 35 -377
rect 41 -381 45 -377
rect 118 -389 122 -385
rect 128 -389 132 -385
rect 151 -389 155 -385
rect 184 -389 188 -385
rect 194 -389 198 -385
rect 736 -357 740 -353
rect 746 -357 750 -353
rect 1146 -357 1150 -353
rect 1156 -357 1160 -353
rect 416 -441 420 -437
rect 430 -441 434 -437
rect 471 -441 475 -437
rect 489 -441 493 -437
rect 524 -441 528 -437
rect 534 -441 538 -437
rect 1248 -441 1252 -437
rect 320 -452 324 -448
rect 330 -452 334 -448
rect 31 -467 35 -463
rect 41 -467 45 -463
rect 119 -505 123 -501
rect 129 -505 133 -501
rect 152 -505 156 -501
rect 185 -505 189 -501
rect 195 -505 199 -501
rect 1262 -441 1266 -437
rect 1303 -441 1307 -437
rect 1321 -441 1325 -437
rect 1356 -441 1360 -437
rect 1366 -441 1370 -437
rect 1146 -452 1150 -448
rect 1156 -452 1160 -448
rect 832 -469 836 -465
rect 846 -469 850 -465
rect 887 -469 891 -465
rect 905 -469 909 -465
rect 940 -469 944 -465
rect 950 -469 954 -465
rect 736 -480 740 -476
rect 746 -480 750 -476
rect 1461 -499 1465 -495
rect 1471 -499 1475 -495
rect 1512 -499 1516 -495
rect 1532 -499 1536 -495
rect 1553 -499 1557 -495
rect 1583 -499 1587 -495
rect 1593 -499 1597 -495
rect 100 -683 104 -679
rect 184 -683 188 -679
rect 231 -683 235 -679
rect 241 -683 245 -679
rect 370 -683 374 -679
rect 454 -683 458 -679
rect 501 -683 505 -679
rect 511 -683 515 -679
<< polysilicon >>
rect 83 60 87 63
rect 104 60 108 63
rect 572 60 576 63
rect 593 60 597 63
rect 956 60 960 63
rect 977 60 981 63
rect 1303 60 1307 63
rect 1324 60 1328 63
rect 83 15 87 52
rect 104 15 108 52
rect 572 15 576 52
rect 593 15 597 52
rect 956 15 960 52
rect 977 15 981 52
rect 1303 15 1307 52
rect 1324 15 1328 52
rect 10 12 14 15
rect 31 12 35 15
rect 499 12 503 15
rect 520 12 524 15
rect 83 4 87 7
rect 10 -33 14 4
rect 31 -33 35 4
rect 104 0 108 7
rect 883 12 887 15
rect 904 12 908 15
rect 572 4 576 7
rect 184 -8 188 -5
rect 205 -8 209 -5
rect 310 -12 314 -9
rect 10 -44 14 -41
rect 31 -49 35 -41
rect 98 -49 102 -46
rect 119 -49 123 -46
rect 184 -53 188 -16
rect 205 -53 209 -16
rect 310 -51 314 -20
rect 499 -33 503 4
rect 520 -33 524 4
rect 593 0 597 7
rect 1230 12 1234 15
rect 1251 12 1255 15
rect 956 4 960 7
rect 673 -8 677 -5
rect 694 -8 698 -5
rect 746 -12 750 -9
rect 499 -44 503 -41
rect 520 -49 524 -41
rect 587 -49 591 -46
rect 608 -49 612 -46
rect 98 -94 102 -57
rect 119 -94 123 -57
rect 673 -53 677 -16
rect 694 -53 698 -16
rect 746 -51 750 -20
rect 883 -33 887 4
rect 904 -33 908 4
rect 977 0 981 7
rect 1303 4 1307 7
rect 1057 -8 1061 -5
rect 1078 -8 1082 -5
rect 1130 -12 1134 -9
rect 883 -44 887 -41
rect 904 -49 908 -41
rect 971 -49 975 -46
rect 992 -49 996 -46
rect 184 -64 188 -61
rect 205 -69 209 -61
rect 310 -62 314 -59
rect 587 -94 591 -57
rect 608 -94 612 -57
rect 1057 -53 1061 -16
rect 1078 -53 1082 -16
rect 1130 -51 1134 -20
rect 1230 -33 1234 4
rect 1251 -33 1255 4
rect 1324 0 1328 7
rect 1404 -8 1408 -5
rect 1425 -8 1429 -5
rect 1477 -12 1481 -9
rect 1230 -44 1234 -41
rect 1251 -49 1255 -41
rect 1318 -49 1322 -46
rect 1339 -49 1343 -46
rect 673 -64 677 -61
rect 694 -69 698 -61
rect 746 -62 750 -59
rect 971 -94 975 -57
rect 992 -94 996 -57
rect 1404 -53 1408 -16
rect 1425 -53 1429 -16
rect 1477 -51 1481 -20
rect 1057 -64 1061 -61
rect 1078 -69 1082 -61
rect 1130 -62 1134 -59
rect 1318 -94 1322 -57
rect 1339 -94 1343 -57
rect 1404 -64 1408 -61
rect 1425 -69 1429 -61
rect 1477 -62 1481 -59
rect 98 -105 102 -102
rect 119 -110 123 -102
rect 587 -105 591 -102
rect 608 -110 612 -102
rect 971 -105 975 -102
rect 992 -110 996 -102
rect 1318 -105 1322 -102
rect 1339 -110 1343 -102
rect 403 -298 407 -295
rect 436 -298 440 -295
rect 460 -298 464 -295
rect 511 -298 515 -295
rect 819 -298 823 -295
rect 852 -298 856 -295
rect 876 -298 880 -295
rect 927 -298 931 -295
rect 1235 -298 1239 -295
rect 1268 -298 1272 -295
rect 1292 -298 1296 -295
rect 1343 -298 1347 -295
rect 325 -351 329 -348
rect 36 -375 40 -372
rect 123 -383 127 -380
rect 144 -383 148 -380
rect 189 -383 193 -380
rect 36 -414 40 -383
rect 36 -425 40 -422
rect 123 -428 127 -391
rect 144 -428 148 -391
rect 189 -428 193 -391
rect 325 -396 329 -359
rect 403 -372 407 -306
rect 436 -372 440 -306
rect 460 -372 464 -306
rect 511 -372 515 -306
rect 741 -351 745 -348
rect 403 -383 407 -380
rect 436 -383 440 -380
rect 460 -383 464 -380
rect 511 -383 515 -380
rect 741 -396 745 -359
rect 819 -372 823 -306
rect 852 -372 856 -306
rect 876 -372 880 -306
rect 927 -372 931 -306
rect 1151 -351 1155 -348
rect 819 -383 823 -380
rect 852 -383 856 -380
rect 876 -383 880 -380
rect 927 -383 931 -380
rect 1151 -396 1155 -359
rect 1235 -372 1239 -306
rect 1268 -372 1272 -306
rect 1292 -372 1296 -306
rect 1343 -372 1347 -306
rect 1235 -383 1239 -380
rect 1268 -383 1272 -380
rect 1292 -383 1296 -380
rect 1343 -383 1347 -380
rect 325 -407 329 -404
rect 741 -407 745 -404
rect 1151 -407 1155 -404
rect 421 -435 425 -432
rect 454 -435 458 -432
rect 478 -435 482 -432
rect 529 -435 533 -432
rect 1253 -435 1257 -432
rect 1286 -435 1290 -432
rect 1310 -435 1314 -432
rect 1361 -435 1365 -432
rect 123 -439 127 -436
rect 144 -444 148 -436
rect 189 -439 193 -436
rect 325 -446 329 -443
rect 36 -461 40 -458
rect 36 -512 40 -469
rect 325 -491 329 -454
rect 124 -499 128 -496
rect 145 -499 149 -496
rect 190 -499 194 -496
rect 325 -502 329 -499
rect 36 -523 40 -520
rect 124 -544 128 -507
rect 145 -544 149 -507
rect 190 -544 194 -507
rect 421 -509 425 -443
rect 454 -509 458 -443
rect 478 -509 482 -443
rect 529 -509 533 -443
rect 1151 -446 1155 -443
rect 837 -463 841 -460
rect 870 -463 874 -460
rect 894 -463 898 -460
rect 945 -463 949 -460
rect 741 -474 745 -471
rect 421 -520 425 -517
rect 454 -520 458 -517
rect 478 -520 482 -517
rect 529 -520 533 -517
rect 741 -519 745 -482
rect 741 -530 745 -527
rect 837 -537 841 -471
rect 870 -537 874 -471
rect 894 -537 898 -471
rect 945 -537 949 -471
rect 1151 -491 1155 -454
rect 1151 -502 1155 -499
rect 1253 -509 1257 -443
rect 1286 -509 1290 -443
rect 1310 -509 1314 -443
rect 1361 -509 1365 -443
rect 1466 -493 1470 -490
rect 1495 -493 1499 -490
rect 1519 -493 1523 -490
rect 1543 -493 1547 -490
rect 1588 -493 1592 -490
rect 1253 -520 1257 -517
rect 1286 -520 1290 -517
rect 1310 -520 1314 -517
rect 1361 -520 1365 -517
rect 1466 -536 1470 -501
rect 1495 -536 1499 -501
rect 1519 -536 1523 -501
rect 1543 -536 1547 -501
rect 1588 -536 1592 -501
rect 837 -548 841 -545
rect 870 -548 874 -545
rect 894 -548 898 -545
rect 945 -548 949 -545
rect 1466 -548 1470 -544
rect 124 -555 128 -552
rect 145 -560 149 -552
rect 190 -555 194 -552
rect 1495 -556 1499 -544
rect 1519 -568 1523 -544
rect 1543 -576 1547 -544
rect 1588 -547 1592 -544
rect 105 -677 109 -674
rect 126 -677 130 -674
rect 147 -677 151 -674
rect 168 -677 172 -674
rect 236 -677 240 -674
rect 375 -677 379 -674
rect 396 -677 400 -674
rect 417 -677 421 -674
rect 438 -677 442 -674
rect 506 -677 510 -674
rect 105 -745 109 -685
rect 126 -745 130 -685
rect 147 -745 151 -685
rect 168 -745 172 -685
rect 236 -745 240 -685
rect 375 -748 379 -685
rect 396 -748 400 -685
rect 417 -748 421 -685
rect 438 -748 442 -685
rect 506 -748 510 -685
rect 105 -756 109 -753
rect 126 -756 130 -753
rect 147 -756 151 -753
rect 168 -756 172 -753
rect 236 -756 240 -753
rect 375 -759 379 -756
rect 396 -759 400 -756
rect 417 -759 421 -756
rect 438 -759 442 -756
rect 506 -759 510 -756
<< polycontact >>
rect 79 33 83 37
rect 568 33 572 37
rect 952 33 956 37
rect 1299 33 1303 37
rect 6 -19 10 -11
rect 100 -1 104 3
rect 180 -35 184 -31
rect 27 -49 31 -45
rect 495 -19 499 -11
rect 306 -39 310 -35
rect 589 -1 593 3
rect 669 -35 673 -31
rect 516 -49 520 -45
rect 94 -76 98 -72
rect 879 -19 883 -11
rect 742 -39 746 -35
rect 973 -1 977 3
rect 1053 -35 1057 -31
rect 900 -49 904 -45
rect 201 -69 205 -65
rect 583 -76 587 -72
rect 1226 -19 1230 -11
rect 1126 -39 1130 -35
rect 1320 -1 1324 3
rect 1400 -35 1404 -31
rect 1247 -49 1251 -45
rect 690 -69 694 -65
rect 967 -76 971 -72
rect 1473 -39 1477 -35
rect 1074 -69 1078 -65
rect 1314 -76 1318 -72
rect 1421 -69 1425 -65
rect 115 -110 119 -106
rect 604 -110 608 -106
rect 988 -110 992 -106
rect 1335 -110 1339 -106
rect 399 -322 403 -318
rect 321 -382 325 -378
rect 32 -402 36 -398
rect 119 -410 123 -406
rect 185 -414 189 -410
rect 432 -330 436 -326
rect 456 -342 460 -338
rect 507 -358 511 -354
rect 815 -322 819 -318
rect 737 -382 741 -378
rect 848 -330 852 -326
rect 872 -342 876 -338
rect 923 -358 927 -354
rect 1231 -322 1235 -318
rect 1147 -382 1151 -378
rect 1264 -330 1268 -326
rect 1288 -342 1292 -338
rect 1339 -358 1343 -354
rect 140 -444 144 -440
rect 32 -500 36 -496
rect 321 -477 325 -473
rect 417 -459 421 -455
rect 120 -526 124 -522
rect 186 -530 190 -526
rect 450 -467 454 -463
rect 474 -479 478 -475
rect 525 -495 529 -491
rect 737 -505 741 -501
rect 833 -487 837 -483
rect 866 -495 870 -491
rect 890 -507 894 -503
rect 941 -523 945 -519
rect 1147 -477 1151 -473
rect 1249 -459 1253 -455
rect 1282 -467 1286 -463
rect 1306 -479 1310 -475
rect 1357 -495 1361 -491
rect 1462 -517 1466 -513
rect 1584 -530 1588 -526
rect 141 -560 145 -556
rect 1491 -556 1495 -552
rect 1515 -568 1519 -564
rect 1539 -576 1543 -572
rect 101 -701 105 -697
rect 122 -709 126 -705
rect 143 -717 147 -713
rect 164 -725 168 -721
rect 232 -733 236 -729
rect 371 -701 375 -697
rect 392 -710 396 -706
rect 413 -719 417 -715
rect 434 -728 438 -724
rect 502 -736 506 -732
<< metal1 >>
rect -202 147 -186 155
rect -170 147 1210 155
rect -202 122 -154 130
rect -138 122 851 130
rect -202 97 -122 105
rect -106 97 479 105
rect -202 72 -87 80
rect -71 72 -49 80
rect 47 76 216 80
rect -65 -11 -49 72
rect -14 60 59 64
rect -14 -11 -10 60
rect 55 37 59 60
rect 78 58 82 76
rect 111 58 115 76
rect 55 33 79 37
rect 88 33 92 54
rect 88 29 156 33
rect 5 25 42 29
rect 5 10 9 25
rect 38 10 42 25
rect 111 13 115 29
rect -65 -19 6 -11
rect 15 -15 19 6
rect 96 -15 100 3
rect 15 -19 100 -15
rect 38 -35 42 -19
rect 23 -107 27 -45
rect 68 -72 72 -19
rect 93 -33 134 -29
rect 152 -31 156 29
rect 179 -10 183 76
rect 212 8 216 76
rect 471 64 479 97
rect 536 76 705 80
rect 471 60 548 64
rect 212 4 309 8
rect 212 -10 216 4
rect 305 -14 309 4
rect 471 -11 479 60
rect 544 37 548 60
rect 567 58 571 76
rect 600 58 604 76
rect 544 33 568 37
rect 577 33 581 54
rect 577 29 645 33
rect 494 25 531 29
rect 494 10 498 25
rect 527 10 531 25
rect 600 13 604 29
rect 93 -51 97 -33
rect 126 -51 130 -33
rect 152 -35 180 -31
rect 189 -35 193 -14
rect 189 -39 306 -35
rect 315 -39 319 -18
rect 471 -19 495 -11
rect 504 -15 508 6
rect 585 -15 589 3
rect 504 -19 589 -15
rect 527 -35 531 -19
rect 212 -55 216 -39
rect 315 -43 351 -39
rect 315 -53 319 -43
rect 68 -76 94 -72
rect 103 -76 107 -55
rect 197 -76 201 -65
rect 103 -80 201 -76
rect 126 -96 130 -80
rect 305 -90 309 -57
rect 512 -72 516 -45
rect 192 -94 309 -90
rect 471 -80 516 -72
rect 557 -72 561 -19
rect 575 -33 623 -29
rect 641 -31 645 29
rect 668 -10 672 76
rect 701 8 705 76
rect 701 4 745 8
rect 701 -10 705 4
rect 741 -14 745 4
rect 843 -11 851 122
rect 920 76 1089 80
rect 859 60 932 64
rect 859 -11 863 60
rect 928 37 932 60
rect 951 58 955 76
rect 984 58 988 76
rect 928 33 952 37
rect 961 33 965 54
rect 961 29 1029 33
rect 878 25 915 29
rect 878 10 882 25
rect 911 10 915 25
rect 984 13 988 29
rect 582 -51 586 -33
rect 615 -51 619 -33
rect 641 -35 669 -31
rect 678 -35 682 -14
rect 678 -39 742 -35
rect 751 -39 755 -18
rect 843 -19 879 -11
rect 888 -15 892 6
rect 969 -15 973 3
rect 888 -19 973 -15
rect 911 -35 915 -19
rect 701 -55 705 -39
rect 751 -43 767 -39
rect 751 -53 755 -43
rect 557 -76 583 -72
rect 592 -76 596 -55
rect 686 -76 690 -65
rect 592 -80 690 -76
rect -202 -115 -55 -107
rect -39 -115 27 -107
rect 23 -125 27 -115
rect 111 -125 115 -106
rect 23 -129 115 -125
rect 162 -124 166 -101
rect 471 -135 479 -80
rect 512 -114 516 -80
rect 615 -96 619 -80
rect 741 -90 745 -57
rect 896 -72 900 -45
rect 681 -94 745 -90
rect 876 -80 900 -72
rect 941 -72 945 -19
rect 959 -33 1007 -29
rect 1025 -31 1029 29
rect 1052 -10 1056 76
rect 1085 8 1089 76
rect 1202 64 1210 147
rect 1267 76 1436 80
rect 1202 60 1279 64
rect 1085 4 1129 8
rect 1085 -10 1089 4
rect 1125 -14 1129 4
rect 1202 -11 1210 60
rect 1275 37 1279 60
rect 1298 58 1302 76
rect 1331 58 1335 76
rect 1275 33 1299 37
rect 1308 33 1312 54
rect 1308 29 1376 33
rect 1225 25 1262 29
rect 1225 10 1229 25
rect 1258 10 1262 25
rect 1331 13 1335 29
rect 966 -51 970 -33
rect 999 -51 1003 -33
rect 1025 -35 1053 -31
rect 1062 -35 1066 -14
rect 1062 -39 1126 -35
rect 1135 -39 1139 -18
rect 1202 -19 1226 -11
rect 1235 -15 1239 6
rect 1316 -15 1320 3
rect 1235 -19 1320 -15
rect 1258 -35 1262 -19
rect 1085 -55 1089 -39
rect 1135 -43 1183 -39
rect 1135 -53 1139 -43
rect 941 -76 967 -72
rect 976 -76 980 -55
rect 1070 -76 1074 -65
rect 976 -80 1074 -76
rect 512 -125 516 -118
rect 600 -125 604 -106
rect 512 -129 604 -125
rect -202 -143 273 -135
rect 289 -143 479 -135
rect 876 -163 884 -80
rect 896 -125 900 -80
rect 999 -96 1003 -80
rect 1125 -90 1129 -57
rect 1243 -72 1247 -45
rect 1065 -94 1129 -90
rect 1198 -80 1247 -72
rect 1288 -72 1292 -19
rect 1306 -33 1354 -29
rect 1372 -31 1376 29
rect 1399 -10 1403 76
rect 1432 8 1436 76
rect 1432 4 1476 8
rect 1432 -10 1436 4
rect 1472 -14 1476 4
rect 1313 -51 1317 -33
rect 1346 -51 1350 -33
rect 1372 -35 1400 -31
rect 1409 -35 1413 -14
rect 1409 -39 1473 -35
rect 1482 -39 1486 -18
rect 1432 -55 1436 -39
rect 1482 -43 1498 -39
rect 1482 -53 1486 -43
rect 1288 -76 1314 -72
rect 1323 -76 1327 -55
rect 1417 -76 1421 -65
rect 1323 -80 1421 -76
rect 984 -125 988 -106
rect 896 -129 988 -125
rect -202 -171 688 -163
rect 704 -171 884 -163
rect 1198 -191 1206 -80
rect 1243 -114 1247 -80
rect 1346 -96 1350 -80
rect 1472 -90 1476 -57
rect 1412 -94 1476 -90
rect 1243 -125 1247 -118
rect 1331 -125 1335 -106
rect 1243 -129 1335 -125
rect -202 -199 1098 -191
rect 1114 -199 1206 -191
rect -101 -215 263 -207
rect -133 -232 682 -224
rect 676 -235 682 -232
rect -144 -257 1092 -249
rect 1086 -260 1092 -257
rect 184 -282 906 -278
rect 911 -282 1465 -278
rect -3 -349 95 -341
rect -3 -369 5 -349
rect -71 -377 5 -369
rect -3 -398 5 -377
rect 31 -359 67 -355
rect 31 -377 35 -359
rect 63 -362 67 -359
rect -3 -402 32 -398
rect 41 -402 45 -381
rect 59 -384 63 -363
rect 59 -388 87 -384
rect 41 -406 75 -402
rect 41 -416 45 -406
rect 31 -430 35 -420
rect 16 -434 35 -430
rect 12 -528 16 -434
rect 31 -445 52 -441
rect 31 -463 35 -445
rect 28 -500 32 -496
rect 41 -500 45 -467
rect 41 -504 53 -500
rect 41 -514 45 -504
rect 31 -528 35 -518
rect 71 -522 75 -406
rect 83 -467 87 -388
rect 91 -419 95 -349
rect 184 -363 188 -282
rect 111 -367 188 -363
rect 118 -385 122 -367
rect 151 -385 155 -367
rect 184 -385 188 -367
rect 263 -318 269 -295
rect 398 -300 402 -282
rect 453 -300 457 -282
rect 506 -300 510 -282
rect 541 -295 545 -282
rect 263 -322 399 -318
rect 263 -378 269 -322
rect 311 -339 324 -335
rect 320 -353 324 -339
rect 263 -382 321 -378
rect 330 -383 334 -357
rect 412 -354 416 -304
rect 471 -354 475 -304
rect 516 -342 520 -304
rect 676 -318 682 -295
rect 814 -300 818 -282
rect 869 -300 873 -282
rect 922 -300 926 -282
rect 676 -322 815 -318
rect 516 -346 580 -342
rect 412 -358 507 -354
rect 471 -374 475 -358
rect 516 -374 520 -346
rect 115 -410 119 -406
rect 128 -410 132 -389
rect 128 -414 185 -410
rect 91 -423 108 -419
rect 104 -452 108 -423
rect 151 -430 155 -414
rect 194 -415 198 -389
rect 330 -387 385 -383
rect 330 -398 334 -387
rect 194 -419 231 -415
rect 320 -415 324 -402
rect 381 -404 385 -387
rect 398 -388 402 -378
rect 506 -388 510 -378
rect 398 -392 514 -388
rect 398 -415 402 -392
rect 541 -415 545 -378
rect 264 -419 402 -415
rect 416 -419 545 -415
rect 194 -430 198 -419
rect 136 -452 140 -440
rect 104 -456 140 -452
rect 83 -471 189 -467
rect 119 -501 123 -471
rect 152 -501 156 -471
rect 185 -501 189 -471
rect 71 -526 120 -522
rect 129 -526 133 -505
rect 12 -532 58 -528
rect 129 -530 186 -526
rect 52 -567 58 -532
rect 105 -568 109 -535
rect 152 -546 156 -530
rect 195 -531 199 -505
rect 195 -535 214 -531
rect 195 -546 199 -535
rect 137 -568 141 -556
rect 105 -572 141 -568
rect 223 -591 231 -419
rect 302 -431 324 -427
rect 298 -537 302 -431
rect 320 -448 324 -431
rect 330 -486 334 -452
rect 330 -490 337 -486
rect 330 -493 334 -490
rect 320 -504 324 -497
rect 345 -504 349 -419
rect 381 -455 385 -428
rect 416 -437 420 -419
rect 471 -437 475 -419
rect 524 -437 528 -419
rect 381 -459 417 -455
rect 430 -491 434 -441
rect 489 -491 493 -441
rect 534 -479 538 -441
rect 534 -483 562 -479
rect 430 -495 525 -491
rect 320 -509 349 -504
rect 489 -511 493 -495
rect 534 -511 538 -483
rect 416 -525 420 -515
rect 524 -525 528 -515
rect 416 -529 528 -525
rect 22 -599 231 -591
rect 268 -541 302 -537
rect 268 -595 279 -541
rect 22 -721 30 -599
rect 572 -607 580 -346
rect 676 -378 682 -322
rect 727 -339 740 -335
rect 736 -353 740 -339
rect 676 -382 737 -378
rect 746 -383 750 -357
rect 828 -354 832 -304
rect 887 -354 891 -304
rect 932 -342 936 -304
rect 1086 -318 1092 -295
rect 1230 -300 1234 -282
rect 1285 -300 1289 -282
rect 1338 -283 1465 -282
rect 1338 -300 1342 -283
rect 1086 -322 1231 -318
rect 932 -346 980 -342
rect 828 -358 923 -354
rect 887 -374 891 -358
rect 932 -374 936 -346
rect 746 -387 801 -383
rect 746 -398 750 -387
rect 736 -443 740 -402
rect 797 -404 801 -387
rect 814 -388 818 -378
rect 922 -388 926 -378
rect 814 -392 926 -388
rect 814 -443 818 -392
rect 922 -419 926 -392
rect 677 -447 818 -443
rect 832 -435 907 -431
rect 718 -459 740 -455
rect 736 -476 740 -459
rect 746 -514 750 -480
rect 746 -518 753 -514
rect 746 -521 750 -518
rect 736 -532 740 -525
rect 761 -532 765 -447
rect 797 -483 801 -456
rect 832 -465 836 -435
rect 887 -465 891 -435
rect 912 -435 944 -431
rect 940 -465 944 -435
rect 797 -487 833 -483
rect 846 -519 850 -469
rect 905 -519 909 -469
rect 950 -507 954 -469
rect 950 -511 962 -507
rect 846 -523 941 -519
rect 736 -533 765 -532
rect 736 -537 820 -533
rect 816 -553 820 -537
rect 905 -539 909 -523
rect 950 -539 954 -511
rect 832 -553 836 -543
rect 940 -553 944 -543
rect 816 -557 944 -553
rect 38 -615 580 -607
rect 38 -713 46 -615
rect 972 -623 980 -346
rect 1086 -378 1092 -322
rect 1137 -339 1150 -335
rect 1146 -353 1150 -339
rect 1086 -382 1147 -378
rect 1156 -383 1160 -357
rect 1244 -354 1248 -304
rect 1303 -354 1307 -304
rect 1348 -342 1352 -304
rect 1348 -346 1396 -342
rect 1244 -358 1339 -354
rect 1303 -374 1307 -358
rect 1348 -374 1352 -346
rect 1156 -387 1217 -383
rect 1156 -398 1160 -387
rect 1146 -415 1150 -402
rect 1213 -404 1217 -387
rect 1230 -388 1234 -378
rect 1338 -388 1342 -378
rect 1230 -392 1342 -388
rect 1230 -415 1234 -392
rect 1087 -419 1234 -415
rect 1248 -419 1360 -415
rect 1088 -525 1092 -419
rect 1128 -431 1150 -427
rect 1146 -448 1150 -431
rect 1156 -486 1160 -452
rect 1156 -490 1163 -486
rect 1156 -493 1160 -490
rect 1146 -504 1150 -497
rect 1171 -504 1175 -419
rect 1213 -455 1217 -428
rect 1248 -437 1252 -419
rect 1303 -437 1307 -419
rect 1356 -437 1360 -419
rect 1213 -459 1249 -455
rect 1262 -491 1266 -441
rect 1321 -491 1325 -441
rect 1366 -479 1370 -441
rect 1366 -483 1378 -479
rect 1262 -495 1357 -491
rect 1146 -509 1175 -504
rect 1321 -511 1325 -495
rect 1366 -511 1370 -483
rect 1248 -525 1252 -515
rect 1356 -525 1360 -515
rect 1088 -529 1360 -525
rect 54 -631 980 -623
rect 54 -705 62 -631
rect 1388 -639 1396 -346
rect 1461 -473 1465 -283
rect 1461 -477 1587 -473
rect 1461 -495 1465 -477
rect 1512 -495 1516 -477
rect 1553 -495 1557 -477
rect 1583 -495 1587 -477
rect 1458 -517 1462 -513
rect 1471 -526 1475 -499
rect 1532 -513 1536 -499
rect 1532 -517 1557 -513
rect 1553 -526 1557 -517
rect 1593 -521 1597 -499
rect 1593 -525 1605 -521
rect 1471 -530 1584 -526
rect 1553 -538 1557 -530
rect 1593 -538 1597 -525
rect 1461 -552 1465 -542
rect 1419 -556 1465 -552
rect 1487 -556 1491 -552
rect 1461 -611 1465 -556
rect 1511 -568 1515 -564
rect 1535 -576 1539 -572
rect 1583 -611 1587 -542
rect 1461 -615 1587 -611
rect 70 -647 1396 -639
rect 70 -697 78 -647
rect 100 -661 505 -657
rect 100 -679 104 -661
rect 231 -679 235 -661
rect 370 -679 374 -661
rect 501 -679 505 -661
rect 70 -701 101 -697
rect 54 -709 122 -705
rect 38 -717 143 -713
rect 22 -725 164 -721
rect 184 -729 188 -683
rect 241 -700 245 -683
rect 241 -704 253 -700
rect 361 -701 371 -697
rect 110 -733 232 -729
rect 110 -747 114 -733
rect 184 -737 188 -733
rect 157 -741 188 -737
rect 157 -747 161 -741
rect 241 -747 245 -704
rect 361 -710 392 -706
rect 361 -719 413 -715
rect 361 -728 434 -724
rect 454 -732 458 -683
rect 511 -714 515 -683
rect 511 -719 522 -714
rect 380 -736 502 -732
rect 380 -750 384 -736
rect 454 -740 458 -736
rect 427 -744 458 -740
rect 427 -750 431 -744
rect 511 -750 515 -719
rect 100 -764 104 -751
rect 133 -764 137 -751
rect 231 -764 235 -751
rect 370 -764 374 -754
rect 403 -764 407 -754
rect 501 -764 505 -754
rect 73 -768 505 -764
<< m2contact >>
rect -186 147 -170 155
rect -154 122 -138 130
rect -122 97 -106 105
rect -87 72 -71 80
rect 42 76 47 81
rect 37 29 42 34
rect 77 4 82 9
rect 4 -44 9 -39
rect 134 -33 139 -28
rect 174 10 179 15
rect 531 76 536 81
rect 526 29 531 34
rect 566 4 571 9
rect 493 -44 498 -39
rect 178 -64 183 -59
rect 187 -94 192 -89
rect 623 -33 628 -28
rect 663 10 668 15
rect 915 76 920 81
rect 910 29 915 34
rect 950 4 955 9
rect 877 -44 882 -39
rect 667 -64 672 -59
rect 92 -105 97 -100
rect 162 -101 167 -96
rect -55 -115 -39 -107
rect 162 -129 170 -124
rect 676 -94 681 -89
rect 1007 -33 1012 -28
rect 1047 10 1052 15
rect 1262 76 1267 81
rect 1257 29 1262 34
rect 1297 4 1302 9
rect 1224 -44 1229 -39
rect 1051 -64 1056 -59
rect 581 -105 586 -100
rect 273 -143 289 -135
rect 1060 -94 1065 -89
rect 1354 -33 1359 -28
rect 1394 10 1399 15
rect 1398 -64 1403 -59
rect 965 -105 970 -100
rect 688 -171 704 -163
rect 1407 -94 1412 -89
rect 1312 -105 1317 -100
rect 1098 -199 1114 -191
rect -106 -215 -101 -207
rect 263 -216 269 -207
rect -138 -232 -133 -224
rect 676 -244 682 -235
rect -149 -257 -144 -249
rect 1086 -269 1092 -260
rect 906 -282 911 -277
rect -87 -377 -71 -369
rect 63 -367 68 -362
rect 11 -434 16 -429
rect 52 -445 57 -440
rect 23 -500 28 -492
rect 53 -504 58 -499
rect 106 -367 111 -362
rect 263 -295 269 -286
rect 306 -287 311 -282
rect 540 -300 545 -295
rect 676 -295 682 -286
rect 722 -287 727 -282
rect 306 -339 311 -334
rect 427 -330 432 -325
rect 1086 -295 1092 -286
rect 1132 -287 1137 -282
rect 540 -378 545 -373
rect 108 -410 115 -405
rect 259 -419 264 -414
rect 514 -392 519 -387
rect 381 -409 386 -404
rect 117 -439 122 -434
rect 183 -439 188 -434
rect 100 -540 105 -535
rect 58 -567 63 -562
rect 214 -535 219 -530
rect 118 -555 123 -550
rect 184 -555 189 -550
rect 297 -431 302 -426
rect 337 -490 342 -485
rect 381 -428 386 -423
rect 445 -467 450 -462
rect 562 -483 567 -478
rect 411 -529 416 -524
rect 268 -600 279 -595
rect 722 -339 727 -334
rect 843 -330 848 -325
rect 1321 -287 1326 -282
rect 672 -447 677 -442
rect 797 -409 802 -404
rect 926 -419 931 -414
rect 713 -459 718 -454
rect 753 -518 758 -513
rect 797 -456 802 -451
rect 907 -436 912 -431
rect 861 -495 866 -490
rect 962 -511 967 -506
rect 1132 -339 1137 -334
rect 1259 -330 1264 -325
rect 1082 -419 1087 -414
rect 1213 -409 1218 -404
rect 1322 -415 1327 -410
rect 1123 -431 1128 -426
rect 1163 -490 1168 -485
rect 1213 -428 1218 -423
rect 1277 -467 1282 -462
rect 1378 -483 1383 -478
rect 1418 -552 1423 -547
rect 268 -657 279 -652
rect 356 -701 361 -696
rect 356 -710 361 -705
rect 356 -719 361 -714
rect 356 -728 361 -723
rect 68 -768 73 -763
<< metal2 >>
rect -186 -249 -170 147
rect -154 -232 -138 122
rect -122 -215 -106 97
rect 38 85 1267 93
rect 38 81 47 85
rect -186 -257 -149 -249
rect -87 -369 -71 72
rect 38 34 42 81
rect 527 81 536 85
rect 527 34 531 81
rect 911 81 920 85
rect 911 34 915 81
rect 1258 81 1267 85
rect 1258 34 1262 81
rect 139 10 174 14
rect 628 10 663 14
rect 1012 10 1047 14
rect 1359 10 1394 14
rect 5 -53 9 -44
rect 78 -53 82 4
rect 139 -28 143 10
rect 139 -33 166 -28
rect -32 -57 82 -53
rect -55 -492 -39 -115
rect -32 -430 -28 -57
rect 78 -114 82 -57
rect 162 -96 166 -33
rect 494 -53 498 -44
rect 567 -53 571 4
rect 628 -33 632 10
rect 494 -57 571 -53
rect 878 -53 882 -44
rect 951 -53 955 4
rect 1012 -33 1016 10
rect 878 -57 955 -53
rect 1225 -53 1229 -44
rect 1298 -53 1302 4
rect 1359 -33 1363 10
rect 1225 -57 1302 -53
rect 179 -90 183 -64
rect 179 -94 187 -90
rect 93 -114 97 -105
rect 179 -114 183 -94
rect 567 -114 571 -57
rect 668 -90 672 -64
rect 668 -94 676 -90
rect 582 -114 586 -105
rect 668 -114 672 -94
rect 951 -114 955 -57
rect 1052 -90 1056 -64
rect 1052 -94 1060 -90
rect 966 -114 970 -105
rect 1052 -114 1056 -94
rect 1298 -114 1302 -57
rect 1399 -90 1403 -64
rect 1399 -94 1407 -90
rect 1313 -114 1317 -105
rect 1399 -114 1403 -94
rect 78 -118 1403 -114
rect 162 -341 170 -129
rect 263 -286 269 -216
rect 107 -349 170 -341
rect 107 -362 111 -349
rect 68 -367 106 -363
rect -32 -434 11 -430
rect 63 -441 69 -367
rect 57 -445 69 -441
rect 77 -410 108 -406
rect -55 -500 23 -492
rect 3 -536 7 -500
rect 77 -500 81 -410
rect 118 -447 122 -439
rect 184 -447 188 -439
rect 255 -447 259 -415
rect 58 -504 81 -500
rect 92 -451 259 -447
rect 92 -527 96 -451
rect 255 -525 259 -451
rect 273 -473 289 -143
rect 307 -334 311 -287
rect 676 -286 682 -244
rect 298 -339 306 -335
rect 371 -330 427 -326
rect 298 -426 302 -339
rect 273 -477 321 -473
rect 311 -513 315 -477
rect 371 -486 375 -330
rect 541 -373 545 -300
rect 519 -392 666 -388
rect 381 -423 385 -409
rect 658 -442 666 -392
rect 658 -447 672 -442
rect 342 -490 375 -486
rect 386 -467 445 -463
rect 386 -513 390 -467
rect 567 -483 596 -479
rect 311 -517 390 -513
rect 92 -531 114 -527
rect 255 -529 411 -525
rect 3 -540 100 -536
rect 110 -563 114 -531
rect 219 -535 247 -531
rect 119 -563 123 -555
rect 185 -563 189 -555
rect 63 -567 189 -563
rect 64 -768 68 -567
rect 239 -582 247 -535
rect 239 -587 314 -582
rect 268 -652 279 -600
rect 306 -724 314 -587
rect 588 -611 596 -483
rect 688 -501 704 -171
rect 723 -334 727 -287
rect 714 -339 722 -335
rect 787 -330 843 -326
rect 714 -454 718 -339
rect 688 -505 737 -501
rect 727 -541 731 -505
rect 787 -514 791 -330
rect 797 -451 801 -409
rect 907 -431 911 -282
rect 1086 -286 1092 -269
rect 931 -419 1082 -414
rect 1098 -473 1114 -199
rect 1133 -334 1137 -287
rect 1124 -339 1132 -335
rect 1203 -330 1259 -326
rect 1124 -426 1128 -339
rect 1098 -477 1147 -473
rect 758 -518 791 -514
rect 802 -495 861 -491
rect 802 -541 806 -495
rect 967 -511 996 -507
rect 727 -545 806 -541
rect 322 -619 596 -611
rect 322 -715 330 -619
rect 988 -627 996 -511
rect 1137 -513 1141 -477
rect 1203 -486 1207 -330
rect 1213 -423 1217 -409
rect 1322 -410 1326 -287
rect 1399 -317 1403 -118
rect 1399 -322 1423 -317
rect 1168 -490 1207 -486
rect 1218 -467 1277 -463
rect 1218 -513 1222 -467
rect 1383 -483 1412 -479
rect 1137 -517 1222 -513
rect 336 -635 996 -627
rect 336 -706 344 -635
rect 1404 -643 1412 -483
rect 1418 -547 1423 -322
rect 348 -651 1412 -643
rect 348 -701 356 -651
rect 336 -710 356 -706
rect 322 -719 356 -715
rect 306 -728 356 -724
<< m123contact >>
rect 351 -43 359 -38
rect 767 -43 775 -37
rect 1183 -43 1191 -38
rect 1498 -43 1506 -37
rect 451 -342 456 -337
rect 469 -479 474 -474
rect 867 -342 872 -337
rect 885 -507 890 -502
rect 1283 -342 1288 -337
rect 1301 -479 1306 -474
rect 1453 -518 1458 -513
rect 1482 -556 1487 -551
rect 1506 -568 1511 -563
rect 1530 -576 1535 -571
<< metal3 >>
rect 351 -338 359 -43
rect 351 -342 451 -338
rect 767 -338 775 -43
rect 767 -342 867 -338
rect 1183 -338 1191 -43
rect 1498 -144 1506 -43
rect 1431 -152 1506 -144
rect 1183 -342 1283 -338
rect 351 -475 359 -342
rect 351 -479 469 -475
rect 351 -595 359 -479
rect 767 -503 775 -342
rect 1183 -475 1191 -342
rect 1183 -479 1301 -475
rect 767 -507 885 -503
rect 767 -583 775 -507
rect 1183 -571 1191 -479
rect 1431 -514 1439 -152
rect 1431 -518 1453 -514
rect 1482 -571 1486 -556
rect 1183 -579 1486 -571
rect 1506 -583 1510 -568
rect 767 -591 1510 -583
rect 1530 -595 1534 -576
rect 351 -603 1534 -595
<< labels >>
rlabel metal1 -200 73 -198 75 3 A3
rlabel metal1 -201 -198 -199 -196 3 B0
rlabel metal2 -2 -497 0 -496 1 B3
rlabel metal1 46 -503 49 -502 1 B3comp
rlabel metal1 48 -405 51 -404 1 A3comp
rlabel metal1 26 -401 29 -400 1 A3
rlabel metal1 -200 -170 -198 -168 3 B1
rlabel metal1 -201 -114 -199 -112 3 B3
rlabel metal2 -31 -56 -28 -54 1 GND
rlabel metal1 -201 -142 -198 -140 2 B2
rlabel metal1 -200 98 -198 100 3 A2
rlabel metal2 46 87 53 91 1 VDD
rlabel metal1 -200 123 -198 125 3 A1
rlabel metal1 -200 149 -198 151 4 A0
rlabel metal1 225 -571 227 -570 1 G3
rlabel metal1 575 -571 578 -570 1 G2
rlabel metal1 974 -571 977 -570 1 G1
rlabel metal3 770 -571 773 -569 1 E2
rlabel metal2 991 -571 994 -570 1 L1
rlabel metal2 732 -504 734 -503 1 B1
rlabel metal2 776 -517 779 -516 1 B1comp
rlabel metal1 958 -510 961 -509 1 L1
rlabel metal1 763 -42 765 -41 1 E2
rlabel metal1 940 -345 943 -344 1 G1
rlabel metal1 754 -386 759 -384 1 A1comp
rlabel metal1 729 -382 734 -380 1 A1
rlabel metal2 591 -571 594 -570 1 L2
rlabel metal1 542 -482 545 -481 1 L2
rlabel metal1 524 -345 527 -344 1 G2
rlabel metal2 242 -571 244 -570 1 L3
rlabel metal1 321 -42 323 -41 1 E3
rlabel metal2 361 -489 363 -488 1 B2comp
rlabel metal1 314 -381 317 -380 1 A2
rlabel metal1 339 -386 342 -385 1 A2comp
rlabel metal2 315 -476 317 -475 1 B2
rlabel metal3 354 -571 357 -569 1 E3
rlabel metal3 1186 -570 1189 -568 1 E1
rlabel metal1 1374 -482 1377 -481 1 L0
rlabel metal1 1356 -345 1359 -344 1 G0
rlabel metal2 1192 -490 1196 -488 1 B0comp
rlabel metal1 1164 -386 1167 -385 1 A0comp
rlabel metal1 1140 -381 1143 -380 1 A0
rlabel metal2 1142 -476 1144 -475 1 B0
rlabel metal1 1390 -570 1393 -568 1 G0
rlabel metal2 1407 -570 1410 -568 1 L0
rlabel metal1 1147 -42 1149 -41 1 E1
rlabel metal1 1493 -42 1495 -41 1 E0
rlabel metal1 1600 -524 1603 -522 7 equal
rlabel metal1 97 -724 99 -723 1 G3
rlabel metal1 97 -716 99 -715 1 G2
rlabel metal1 97 -708 99 -707 1 G1
rlabel metal1 97 -700 99 -699 1 G0
rlabel metal1 246 -703 248 -702 1 greater
rlabel metal1 364 -700 366 -699 1 L0
rlabel metal1 364 -709 366 -708 1 L1
rlabel metal1 364 -718 366 -717 1 L2
rlabel metal1 364 -727 366 -726 1 L3
rlabel metal1 517 -718 519 -717 1 lesser
<< end >>
