* SPICE3 file created from not.ext - technology: scmos
.include TSMC_180nm.txt

.param SUPPLY = 1.8
.param LAMBDA = 0.18u
.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}
.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd VDD gnd 'Supply'

Vin_not Vin gnd DC(0)

.option scale=0.09u

M1000 Vout Vin GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=48 ps=28
M1001 Vout Vin VDD w_n2_0# CMOSP w=8 l=4
+  ad=48 pd=28 as=48 ps=28
C0 Vin Vout 0.03fF
C1 Vout w_n2_0# 0.03fF
C2 VDD Vout 0.03fF
C3 Vin w_n2_0# 0.11fF
C4 Vout GND 0.03fF
C5 VDD w_n2_0# 0.03fF
C6 GND Gnd 0.08fF
C7 Vout Gnd 0.08fF
C8 VDD Gnd 0.08fF
C9 Vin Gnd 0.27fF
C10 w_n2_0# Gnd 0.67fF

.tran 1n 800n

.control
run
plot v(Vout)+2 v(Vin)

.end
.endc
