magic
tech scmos
timestamp 1700524057
<< nwell >>
rect 148 782 208 806
rect 214 782 242 806
rect 145 690 205 714
rect 211 690 239 714
rect 145 598 205 622
rect 211 598 239 622
rect 145 506 205 530
rect 211 506 239 530
rect 150 415 210 439
rect 216 415 244 439
rect 147 323 207 347
rect 213 323 241 347
rect 147 231 207 255
rect 213 231 241 255
rect 147 139 207 163
rect 213 139 241 163
<< ntransistor >>
rect 160 745 164 753
rect 181 745 185 753
rect 226 745 230 753
rect 157 653 161 661
rect 178 653 182 661
rect 223 653 227 661
rect 157 561 161 569
rect 178 561 182 569
rect 223 561 227 569
rect 157 469 161 477
rect 178 469 182 477
rect 223 469 227 477
rect 162 378 166 386
rect 183 378 187 386
rect 228 378 232 386
rect 159 286 163 294
rect 180 286 184 294
rect 225 286 229 294
rect 159 194 163 202
rect 180 194 184 202
rect 225 194 229 202
rect 159 102 163 110
rect 180 102 184 110
rect 225 102 229 110
<< ptransistor >>
rect 160 790 164 798
rect 181 790 185 798
rect 226 790 230 798
rect 157 698 161 706
rect 178 698 182 706
rect 223 698 227 706
rect 157 606 161 614
rect 178 606 182 614
rect 223 606 227 614
rect 157 514 161 522
rect 178 514 182 522
rect 223 514 227 522
rect 162 423 166 431
rect 183 423 187 431
rect 228 423 232 431
rect 159 331 163 339
rect 180 331 184 339
rect 225 331 229 339
rect 159 239 163 247
rect 180 239 184 247
rect 225 239 229 247
rect 159 147 163 155
rect 180 147 184 155
rect 225 147 229 155
<< ndiffusion >>
rect 154 751 160 753
rect 154 747 155 751
rect 159 747 160 751
rect 154 745 160 747
rect 164 745 181 753
rect 185 751 202 753
rect 185 747 188 751
rect 192 747 202 751
rect 185 745 202 747
rect 220 751 226 753
rect 220 747 221 751
rect 225 747 226 751
rect 220 745 226 747
rect 230 751 236 753
rect 230 747 231 751
rect 235 747 236 751
rect 230 745 236 747
rect 151 659 157 661
rect 151 655 152 659
rect 156 655 157 659
rect 151 653 157 655
rect 161 653 178 661
rect 182 659 199 661
rect 182 655 185 659
rect 189 655 199 659
rect 182 653 199 655
rect 217 659 223 661
rect 217 655 218 659
rect 222 655 223 659
rect 217 653 223 655
rect 227 659 233 661
rect 227 655 228 659
rect 232 655 233 659
rect 227 653 233 655
rect 151 567 157 569
rect 151 563 152 567
rect 156 563 157 567
rect 151 561 157 563
rect 161 561 178 569
rect 182 567 199 569
rect 182 563 185 567
rect 189 563 199 567
rect 182 561 199 563
rect 217 567 223 569
rect 217 563 218 567
rect 222 563 223 567
rect 217 561 223 563
rect 227 567 233 569
rect 227 563 228 567
rect 232 563 233 567
rect 227 561 233 563
rect 151 475 157 477
rect 151 471 152 475
rect 156 471 157 475
rect 151 469 157 471
rect 161 469 178 477
rect 182 475 199 477
rect 182 471 185 475
rect 189 471 199 475
rect 182 469 199 471
rect 217 475 223 477
rect 217 471 218 475
rect 222 471 223 475
rect 217 469 223 471
rect 227 475 233 477
rect 227 471 228 475
rect 232 471 233 475
rect 227 469 233 471
rect 156 384 162 386
rect 156 380 157 384
rect 161 380 162 384
rect 156 378 162 380
rect 166 378 183 386
rect 187 384 204 386
rect 187 380 190 384
rect 194 380 204 384
rect 187 378 204 380
rect 222 384 228 386
rect 222 380 223 384
rect 227 380 228 384
rect 222 378 228 380
rect 232 384 238 386
rect 232 380 233 384
rect 237 380 238 384
rect 232 378 238 380
rect 153 292 159 294
rect 153 288 154 292
rect 158 288 159 292
rect 153 286 159 288
rect 163 286 180 294
rect 184 292 201 294
rect 184 288 187 292
rect 191 288 201 292
rect 184 286 201 288
rect 219 292 225 294
rect 219 288 220 292
rect 224 288 225 292
rect 219 286 225 288
rect 229 292 235 294
rect 229 288 230 292
rect 234 288 235 292
rect 229 286 235 288
rect 153 200 159 202
rect 153 196 154 200
rect 158 196 159 200
rect 153 194 159 196
rect 163 194 180 202
rect 184 200 201 202
rect 184 196 187 200
rect 191 196 201 200
rect 184 194 201 196
rect 219 200 225 202
rect 219 196 220 200
rect 224 196 225 200
rect 219 194 225 196
rect 229 200 235 202
rect 229 196 230 200
rect 234 196 235 200
rect 229 194 235 196
rect 153 108 159 110
rect 153 104 154 108
rect 158 104 159 108
rect 153 102 159 104
rect 163 102 180 110
rect 184 108 201 110
rect 184 104 187 108
rect 191 104 201 108
rect 184 102 201 104
rect 219 108 225 110
rect 219 104 220 108
rect 224 104 225 108
rect 219 102 225 104
rect 229 108 235 110
rect 229 104 230 108
rect 234 104 235 108
rect 229 102 235 104
<< pdiffusion >>
rect 154 796 160 798
rect 154 792 155 796
rect 159 792 160 796
rect 154 790 160 792
rect 164 796 181 798
rect 164 792 165 796
rect 169 792 181 796
rect 164 790 181 792
rect 185 796 202 798
rect 185 792 188 796
rect 192 792 202 796
rect 185 790 202 792
rect 220 796 226 798
rect 220 792 221 796
rect 225 792 226 796
rect 220 790 226 792
rect 230 796 236 798
rect 230 792 231 796
rect 235 792 236 796
rect 230 790 236 792
rect 151 704 157 706
rect 151 700 152 704
rect 156 700 157 704
rect 151 698 157 700
rect 161 704 178 706
rect 161 700 162 704
rect 166 700 178 704
rect 161 698 178 700
rect 182 704 199 706
rect 182 700 185 704
rect 189 700 199 704
rect 182 698 199 700
rect 217 704 223 706
rect 217 700 218 704
rect 222 700 223 704
rect 217 698 223 700
rect 227 704 233 706
rect 227 700 228 704
rect 232 700 233 704
rect 227 698 233 700
rect 151 612 157 614
rect 151 608 152 612
rect 156 608 157 612
rect 151 606 157 608
rect 161 612 178 614
rect 161 608 162 612
rect 166 608 178 612
rect 161 606 178 608
rect 182 612 199 614
rect 182 608 185 612
rect 189 608 199 612
rect 182 606 199 608
rect 217 612 223 614
rect 217 608 218 612
rect 222 608 223 612
rect 217 606 223 608
rect 227 612 233 614
rect 227 608 228 612
rect 232 608 233 612
rect 227 606 233 608
rect 151 520 157 522
rect 151 516 152 520
rect 156 516 157 520
rect 151 514 157 516
rect 161 520 178 522
rect 161 516 162 520
rect 166 516 178 520
rect 161 514 178 516
rect 182 520 199 522
rect 182 516 185 520
rect 189 516 199 520
rect 182 514 199 516
rect 217 520 223 522
rect 217 516 218 520
rect 222 516 223 520
rect 217 514 223 516
rect 227 520 233 522
rect 227 516 228 520
rect 232 516 233 520
rect 227 514 233 516
rect 156 429 162 431
rect 156 425 157 429
rect 161 425 162 429
rect 156 423 162 425
rect 166 429 183 431
rect 166 425 167 429
rect 171 425 183 429
rect 166 423 183 425
rect 187 429 204 431
rect 187 425 190 429
rect 194 425 204 429
rect 187 423 204 425
rect 222 429 228 431
rect 222 425 223 429
rect 227 425 228 429
rect 222 423 228 425
rect 232 429 238 431
rect 232 425 233 429
rect 237 425 238 429
rect 232 423 238 425
rect 153 337 159 339
rect 153 333 154 337
rect 158 333 159 337
rect 153 331 159 333
rect 163 337 180 339
rect 163 333 164 337
rect 168 333 180 337
rect 163 331 180 333
rect 184 337 201 339
rect 184 333 187 337
rect 191 333 201 337
rect 184 331 201 333
rect 219 337 225 339
rect 219 333 220 337
rect 224 333 225 337
rect 219 331 225 333
rect 229 337 235 339
rect 229 333 230 337
rect 234 333 235 337
rect 229 331 235 333
rect 153 245 159 247
rect 153 241 154 245
rect 158 241 159 245
rect 153 239 159 241
rect 163 245 180 247
rect 163 241 164 245
rect 168 241 180 245
rect 163 239 180 241
rect 184 245 201 247
rect 184 241 187 245
rect 191 241 201 245
rect 184 239 201 241
rect 219 245 225 247
rect 219 241 220 245
rect 224 241 225 245
rect 219 239 225 241
rect 229 245 235 247
rect 229 241 230 245
rect 234 241 235 245
rect 229 239 235 241
rect 153 153 159 155
rect 153 149 154 153
rect 158 149 159 153
rect 153 147 159 149
rect 163 153 180 155
rect 163 149 164 153
rect 168 149 180 153
rect 163 147 180 149
rect 184 153 201 155
rect 184 149 187 153
rect 191 149 201 153
rect 184 147 201 149
rect 219 153 225 155
rect 219 149 220 153
rect 224 149 225 153
rect 219 147 225 149
rect 229 153 235 155
rect 229 149 230 153
rect 234 149 235 153
rect 229 147 235 149
<< ndcontact >>
rect 155 747 159 751
rect 188 747 192 751
rect 221 747 225 751
rect 231 747 235 751
rect 152 655 156 659
rect 185 655 189 659
rect 218 655 222 659
rect 228 655 232 659
rect 152 563 156 567
rect 185 563 189 567
rect 218 563 222 567
rect 228 563 232 567
rect 152 471 156 475
rect 185 471 189 475
rect 218 471 222 475
rect 228 471 232 475
rect 157 380 161 384
rect 190 380 194 384
rect 223 380 227 384
rect 233 380 237 384
rect 154 288 158 292
rect 187 288 191 292
rect 220 288 224 292
rect 230 288 234 292
rect 154 196 158 200
rect 187 196 191 200
rect 220 196 224 200
rect 230 196 234 200
rect 154 104 158 108
rect 187 104 191 108
rect 220 104 224 108
rect 230 104 234 108
<< pdcontact >>
rect 155 792 159 796
rect 165 792 169 796
rect 188 792 192 796
rect 221 792 225 796
rect 231 792 235 796
rect 152 700 156 704
rect 162 700 166 704
rect 185 700 189 704
rect 218 700 222 704
rect 228 700 232 704
rect 152 608 156 612
rect 162 608 166 612
rect 185 608 189 612
rect 218 608 222 612
rect 228 608 232 612
rect 152 516 156 520
rect 162 516 166 520
rect 185 516 189 520
rect 218 516 222 520
rect 228 516 232 520
rect 157 425 161 429
rect 167 425 171 429
rect 190 425 194 429
rect 223 425 227 429
rect 233 425 237 429
rect 154 333 158 337
rect 164 333 168 337
rect 187 333 191 337
rect 220 333 224 337
rect 230 333 234 337
rect 154 241 158 245
rect 164 241 168 245
rect 187 241 191 245
rect 220 241 224 245
rect 230 241 234 245
rect 154 149 158 153
rect 164 149 168 153
rect 187 149 191 153
rect 220 149 224 153
rect 230 149 234 153
<< polysilicon >>
rect 160 798 164 801
rect 181 798 185 801
rect 226 798 230 801
rect 160 753 164 790
rect 181 753 185 790
rect 226 753 230 790
rect 160 742 164 745
rect 181 742 185 745
rect 226 742 230 745
rect 157 706 161 709
rect 178 706 182 709
rect 223 706 227 709
rect 157 661 161 698
rect 178 661 182 698
rect 223 661 227 698
rect 157 650 161 653
rect 178 650 182 653
rect 223 650 227 653
rect 157 614 161 617
rect 178 614 182 617
rect 223 614 227 617
rect 157 569 161 606
rect 178 569 182 606
rect 223 569 227 606
rect 157 558 161 561
rect 178 558 182 561
rect 223 558 227 561
rect 157 522 161 525
rect 178 522 182 525
rect 223 522 227 525
rect 157 477 161 514
rect 178 477 182 514
rect 223 477 227 514
rect 157 466 161 469
rect 178 466 182 469
rect 223 466 227 469
rect 162 431 166 434
rect 183 431 187 434
rect 228 431 232 434
rect 162 386 166 423
rect 183 386 187 423
rect 228 386 232 423
rect 162 375 166 378
rect 183 375 187 378
rect 228 375 232 378
rect 159 339 163 342
rect 180 339 184 342
rect 225 339 229 342
rect 159 294 163 331
rect 180 294 184 331
rect 225 294 229 331
rect 159 283 163 286
rect 180 283 184 286
rect 225 283 229 286
rect 159 247 163 250
rect 180 247 184 250
rect 225 247 229 250
rect 159 202 163 239
rect 180 202 184 239
rect 225 202 229 239
rect 159 191 163 194
rect 180 191 184 194
rect 225 191 229 194
rect 159 155 163 158
rect 180 155 184 158
rect 225 155 229 158
rect 159 110 163 147
rect 180 110 184 147
rect 225 110 229 147
rect 159 99 163 102
rect 180 99 184 102
rect 225 99 229 102
<< polycontact >>
rect 156 771 160 775
rect 177 759 181 763
rect 222 767 226 771
rect 153 679 157 683
rect 174 667 178 671
rect 219 675 223 679
rect 153 587 157 591
rect 174 575 178 579
rect 219 583 223 587
rect 153 495 157 499
rect 174 483 178 487
rect 219 491 223 495
rect 158 404 162 408
rect 179 392 183 396
rect 224 400 228 404
rect 155 312 159 316
rect 176 300 180 304
rect 221 308 225 312
rect 155 220 159 224
rect 176 208 180 212
rect 221 216 225 220
rect 155 128 159 132
rect 176 116 180 120
rect 221 124 225 128
<< metal1 >>
rect 126 763 130 826
rect 146 814 225 818
rect 155 796 159 814
rect 188 796 192 814
rect 221 796 225 814
rect 146 771 156 775
rect 165 771 169 792
rect 165 767 222 771
rect 126 759 177 763
rect 126 671 130 759
rect 188 751 192 767
rect 231 766 235 792
rect 231 762 242 766
rect 231 751 235 762
rect 155 737 159 747
rect 221 737 225 747
rect 155 733 225 737
rect 146 723 222 727
rect 152 704 156 723
rect 185 704 189 723
rect 218 704 222 723
rect 146 679 153 683
rect 162 679 166 700
rect 162 675 219 679
rect 126 667 174 671
rect 126 579 130 667
rect 185 659 189 675
rect 228 674 232 700
rect 228 670 239 674
rect 228 659 232 670
rect 152 645 156 655
rect 218 645 222 655
rect 152 641 222 645
rect 146 631 222 635
rect 152 612 156 631
rect 185 612 189 631
rect 218 612 222 631
rect 146 587 153 591
rect 162 587 166 608
rect 162 583 219 587
rect 126 575 174 579
rect 126 487 130 575
rect 185 567 189 583
rect 228 582 232 608
rect 228 578 239 582
rect 228 567 232 578
rect 152 553 156 563
rect 218 553 222 563
rect 152 549 222 553
rect 146 539 222 543
rect 152 520 156 539
rect 185 520 189 539
rect 218 520 222 539
rect 146 495 153 499
rect 162 495 166 516
rect 162 491 219 495
rect 126 483 174 487
rect 126 396 130 483
rect 185 475 189 491
rect 228 490 232 516
rect 228 486 239 490
rect 228 475 232 486
rect 152 461 156 471
rect 218 461 222 471
rect 152 457 222 461
rect 148 447 227 451
rect 157 429 161 447
rect 190 429 194 447
rect 223 429 227 447
rect 148 404 158 408
rect 167 404 171 425
rect 167 400 224 404
rect 126 392 179 396
rect 126 304 130 392
rect 190 384 194 400
rect 233 399 237 425
rect 233 395 241 399
rect 233 384 237 395
rect 157 370 161 380
rect 223 370 227 380
rect 157 366 227 370
rect 148 356 224 360
rect 154 337 158 356
rect 187 337 191 356
rect 220 337 224 356
rect 148 312 155 316
rect 164 312 168 333
rect 164 308 221 312
rect 126 300 176 304
rect 126 212 130 300
rect 187 292 191 308
rect 230 307 234 333
rect 230 303 241 307
rect 230 292 234 303
rect 154 278 158 288
rect 220 278 224 288
rect 154 274 224 278
rect 148 264 224 268
rect 154 245 158 264
rect 187 245 191 264
rect 220 245 224 264
rect 148 220 155 224
rect 164 220 168 241
rect 164 216 221 220
rect 126 208 176 212
rect 126 120 130 208
rect 187 200 191 216
rect 230 215 234 241
rect 230 211 241 215
rect 230 200 234 211
rect 154 186 158 196
rect 220 186 224 196
rect 154 182 224 186
rect 148 172 224 176
rect 154 153 158 172
rect 187 153 191 172
rect 220 153 224 172
rect 148 128 155 132
rect 164 128 168 149
rect 164 124 221 128
rect 126 116 176 120
rect 187 108 191 124
rect 230 123 234 149
rect 230 119 241 123
rect 230 108 234 119
rect 154 94 158 104
rect 220 94 224 104
rect 154 90 224 94
<< m2contact >>
rect 141 771 146 776
rect 225 733 230 738
rect 141 679 146 684
rect 222 641 227 646
rect 141 587 146 592
rect 222 549 227 554
rect 141 495 146 500
rect 222 457 227 462
rect 143 404 148 409
rect 227 366 232 371
rect 143 312 148 317
rect 224 274 229 279
rect 143 220 148 225
rect 224 182 229 187
rect 143 128 148 133
rect 224 90 229 95
<< metal2 >>
rect 110 771 141 775
rect 248 737 252 826
rect 230 733 252 737
rect 110 679 141 683
rect 248 645 252 733
rect 227 641 252 645
rect 110 587 141 591
rect 248 553 252 641
rect 227 549 252 553
rect 110 495 141 499
rect 248 461 252 549
rect 227 457 252 461
rect 110 404 143 408
rect 248 370 252 457
rect 232 366 252 370
rect 110 312 143 316
rect 248 278 252 366
rect 229 274 252 278
rect 110 220 143 224
rect 248 186 252 274
rect 229 182 252 186
rect 110 128 143 132
rect 248 94 252 182
rect 229 90 252 94
<< m123contact >>
rect 141 814 146 819
rect 141 723 146 728
rect 141 631 146 636
rect 141 539 146 544
rect 143 447 148 452
rect 143 356 148 361
rect 143 264 148 269
rect 143 172 148 177
<< metal3 >>
rect 118 814 141 818
rect 118 727 122 814
rect 118 723 141 727
rect 118 635 122 723
rect 118 631 141 635
rect 118 543 122 631
rect 118 539 141 543
rect 118 451 122 539
rect 118 447 143 451
rect 118 360 122 447
rect 118 356 143 360
rect 118 268 122 356
rect 118 264 143 268
rect 118 176 122 264
rect 118 172 143 176
<< labels >>
rlabel metal2 112 772 115 774 3 A3
rlabel metal3 119 814 122 816 5 VDD
rlabel metal1 236 764 239 765 1 A3out
rlabel metal2 111 681 114 683 3 A2
rlabel metal1 233 671 236 672 1 A2out
rlabel metal2 113 589 116 591 3 A1
rlabel metal1 233 579 236 580 1 A1out
rlabel metal2 111 495 114 497 3 A0
rlabel metal1 234 487 237 488 1 A0out
rlabel metal2 112 406 115 408 3 B3
rlabel metal1 236 304 239 305 1 B2out
rlabel metal2 112 313 115 315 3 B2
rlabel metal2 111 221 113 222 3 B1
rlabel metal1 235 212 238 213 1 B1out
rlabel metal2 111 129 114 130 3 B0
rlabel metal1 236 120 239 121 1 B0out
rlabel metal1 236 396 239 397 1 B3out
rlabel metal2 250 822 252 824 6 GND
rlabel metal1 126 822 128 823 5 E
<< end >>
