magic
tech scmos
timestamp 1700489452
<< nwell >>
rect -2 0 91 24
rect 99 0 127 24
<< ntransistor >>
rect 10 -44 14 -36
rect 39 -44 43 -36
rect 63 -44 67 -36
rect 111 -44 115 -36
<< ptransistor >>
rect 10 8 14 16
rect 39 8 43 16
rect 63 8 67 16
rect 111 8 115 16
<< ndiffusion >>
rect 4 -38 10 -36
rect 4 -42 5 -38
rect 9 -42 10 -38
rect 4 -44 10 -42
rect 14 -44 39 -36
rect 43 -44 63 -36
rect 67 -38 85 -36
rect 67 -42 74 -38
rect 78 -42 85 -38
rect 67 -44 85 -42
rect 105 -38 111 -36
rect 105 -42 106 -38
rect 110 -42 111 -38
rect 105 -44 111 -42
rect 115 -38 121 -36
rect 115 -42 116 -38
rect 120 -42 121 -38
rect 115 -44 121 -42
<< pdiffusion >>
rect 4 14 10 16
rect 4 10 5 14
rect 9 10 10 14
rect 4 8 10 10
rect 14 14 39 16
rect 14 10 15 14
rect 19 10 39 14
rect 14 8 39 10
rect 43 14 63 16
rect 43 10 56 14
rect 60 10 63 14
rect 43 8 63 10
rect 67 14 85 16
rect 67 10 74 14
rect 78 10 85 14
rect 67 8 85 10
rect 105 14 111 16
rect 105 10 106 14
rect 110 10 111 14
rect 105 8 111 10
rect 115 14 121 16
rect 115 10 116 14
rect 120 10 121 14
rect 115 8 121 10
<< ndcontact >>
rect 5 -42 9 -38
rect 74 -42 78 -38
rect 106 -42 110 -38
rect 116 -42 120 -38
<< pdcontact >>
rect 5 10 9 14
rect 15 10 19 14
rect 56 10 60 14
rect 74 10 78 14
rect 106 10 110 14
rect 116 10 120 14
<< polysilicon >>
rect 10 16 14 19
rect 39 16 43 19
rect 63 16 67 19
rect 111 16 115 19
rect 10 -36 14 8
rect 39 -36 43 8
rect 63 -36 67 8
rect 111 -36 115 8
rect 10 -47 14 -44
rect 39 -47 43 -44
rect 63 -47 67 -44
rect 111 -47 115 -44
<< polycontact >>
rect 6 -8 10 -4
rect 35 -24 39 -20
rect 59 -32 63 -28
rect 107 -16 111 -12
<< metal1 >>
rect -2 32 127 36
rect 5 14 9 32
rect 56 14 60 32
rect 106 14 110 32
rect 2 -8 6 -4
rect 15 -12 19 10
rect 74 -12 78 10
rect 15 -16 107 -12
rect 2 -24 35 -20
rect 2 -32 59 -28
rect 74 -38 78 -16
rect 116 -20 120 10
rect 116 -24 128 -20
rect 116 -38 120 -24
rect 5 -52 9 -42
rect 106 -52 110 -42
rect -2 -56 119 -52
<< labels >>
rlabel metal1 2 34 4 35 4 VDD
rlabel metal1 3 -7 5 -6 1 VA
rlabel metal1 2 -55 4 -54 2 GND
rlabel metal1 123 -23 125 -22 7 Vout
rlabel metal1 3 -23 5 -22 1 VB
rlabel metal1 3 -31 5 -30 1 VC
<< end >>
