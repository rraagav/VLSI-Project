magic
tech scmos
timestamp 1700488278
<< nwell >>
rect -2 0 58 24
rect 64 0 92 24
<< ntransistor >>
rect 10 -37 14 -29
rect 31 -37 35 -29
rect 76 -37 80 -29
<< ptransistor >>
rect 10 8 14 16
rect 31 8 35 16
rect 76 8 80 16
<< ndiffusion >>
rect 4 -31 10 -29
rect 4 -35 5 -31
rect 9 -35 10 -31
rect 4 -37 10 -35
rect 14 -37 31 -29
rect 35 -31 52 -29
rect 35 -35 38 -31
rect 42 -35 52 -31
rect 35 -37 52 -35
rect 70 -31 76 -29
rect 70 -35 71 -31
rect 75 -35 76 -31
rect 70 -37 76 -35
rect 80 -31 86 -29
rect 80 -35 81 -31
rect 85 -35 86 -31
rect 80 -37 86 -35
<< pdiffusion >>
rect 4 14 10 16
rect 4 10 5 14
rect 9 10 10 14
rect 4 8 10 10
rect 14 14 31 16
rect 14 10 15 14
rect 19 10 31 14
rect 14 8 31 10
rect 35 14 52 16
rect 35 10 38 14
rect 42 10 52 14
rect 35 8 52 10
rect 70 14 76 16
rect 70 10 71 14
rect 75 10 76 14
rect 70 8 76 10
rect 80 14 86 16
rect 80 10 81 14
rect 85 10 86 14
rect 80 8 86 10
<< ndcontact >>
rect 5 -35 9 -31
rect 38 -35 42 -31
rect 71 -35 75 -31
rect 81 -35 85 -31
<< pdcontact >>
rect 5 10 9 14
rect 15 10 19 14
rect 38 10 42 14
rect 71 10 75 14
rect 81 10 85 14
<< polysilicon >>
rect 10 16 14 19
rect 31 16 35 19
rect 76 16 80 19
rect 10 -29 14 8
rect 31 -29 35 8
rect 76 -29 80 8
rect 10 -40 14 -37
rect 31 -40 35 -37
rect 76 -40 80 -37
<< polycontact >>
rect 6 -11 10 -7
rect 27 -23 31 -19
rect 72 -15 76 -11
<< metal1 >>
rect -2 32 75 36
rect 5 14 9 32
rect 38 14 42 32
rect 71 14 75 32
rect 2 -11 6 -7
rect 15 -11 19 10
rect 15 -15 72 -11
rect 2 -23 27 -19
rect 38 -31 42 -15
rect 81 -16 85 10
rect 81 -20 92 -16
rect 81 -31 85 -20
rect 5 -45 9 -35
rect 71 -45 75 -35
rect -2 -49 75 -45
<< labels >>
rlabel metal1 86 -19 88 -18 7 Vout
rlabel metal1 2 34 4 35 4 VDD
rlabel metal1 2 -48 4 -47 2 GND
rlabel metal1 3 -10 5 -9 1 VA
rlabel metal1 3 -22 5 -21 1 VB
<< end >>
