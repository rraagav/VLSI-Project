magic
tech scmos
timestamp 1700544712
<< nwell >>
rect -884 131 -856 155
rect -808 131 -748 155
rect -742 131 -714 155
rect -638 131 -578 155
rect -572 131 -544 155
rect -881 22 -853 46
rect -808 22 -748 46
rect -742 22 -714 46
rect -642 22 -582 46
rect -576 22 -548 46
rect -448 22 -420 46
rect -159 -32 -99 -8
rect 439 -32 499 -8
rect 1318 -32 1378 -8
rect 2086 -32 2146 -8
rect -232 -80 -172 -56
rect -58 -100 2 -76
rect 366 -80 426 -56
rect 540 -100 600 -76
rect 1245 -80 1305 -56
rect 1419 -100 1479 -76
rect 2013 -80 2073 -56
rect 2187 -100 2247 -76
rect -586 -133 -526 -109
rect -520 -133 -492 -109
rect -144 -141 -84 -117
rect 454 -141 514 -117
rect 1333 -141 1393 -117
rect 2101 -141 2161 -117
rect -589 -225 -529 -201
rect -523 -225 -495 -201
rect -589 -317 -529 -293
rect -523 -317 -495 -293
rect 122 -335 182 -311
rect 865 -338 925 -314
rect 1624 -338 1684 -314
rect 2360 -338 2420 -314
rect -188 -383 -128 -359
rect 49 -383 109 -359
rect -589 -409 -529 -385
rect -523 -409 -495 -385
rect 223 -403 283 -379
rect 555 -386 615 -362
rect 792 -386 852 -362
rect 966 -406 1026 -382
rect 1314 -386 1374 -362
rect 1551 -386 1611 -362
rect 1725 -406 1785 -382
rect 2050 -386 2110 -362
rect 2287 -386 2347 -362
rect 2461 -406 2521 -382
rect -261 -431 -201 -407
rect -87 -451 -27 -427
rect 137 -444 197 -420
rect 482 -434 542 -410
rect 656 -454 716 -430
rect 880 -447 940 -423
rect 1241 -434 1301 -410
rect 1415 -454 1475 -430
rect 1639 -447 1699 -423
rect 1977 -434 2037 -410
rect 2151 -454 2211 -430
rect 2375 -447 2435 -423
rect -584 -500 -524 -476
rect -518 -500 -490 -476
rect -173 -492 -113 -468
rect 570 -495 630 -471
rect 1329 -495 1389 -471
rect 2065 -495 2125 -471
rect 109 -550 169 -526
rect 175 -550 203 -526
rect 268 -550 328 -526
rect 336 -550 364 -526
rect 852 -553 912 -529
rect 918 -553 946 -529
rect 1011 -553 1071 -529
rect 1079 -553 1107 -529
rect 1611 -553 1671 -529
rect 1677 -553 1705 -529
rect 1770 -553 1830 -529
rect 1838 -553 1866 -529
rect 2347 -553 2407 -529
rect 2413 -553 2441 -529
rect 2506 -553 2566 -529
rect 2574 -553 2602 -529
rect -587 -592 -527 -568
rect -521 -592 -493 -568
rect -202 -601 -142 -577
rect -136 -601 -108 -577
rect 541 -604 601 -580
rect 607 -604 635 -580
rect 1300 -604 1360 -580
rect 1366 -604 1394 -580
rect 2036 -604 2096 -580
rect 2102 -604 2130 -580
rect -587 -684 -527 -660
rect -521 -684 -493 -660
rect -587 -776 -527 -752
rect -521 -776 -493 -752
rect -130 -825 -70 -801
rect 468 -825 528 -801
rect 1347 -825 1407 -801
rect 2115 -825 2175 -801
rect -203 -873 -143 -849
rect -29 -893 31 -869
rect 395 -873 455 -849
rect 569 -893 629 -869
rect 1274 -873 1334 -849
rect 1448 -893 1508 -869
rect 2042 -873 2102 -849
rect 2216 -893 2276 -869
rect -586 -926 -526 -902
rect -520 -926 -492 -902
rect -115 -934 -55 -910
rect 483 -934 543 -910
rect 1362 -934 1422 -910
rect 2130 -934 2190 -910
rect -589 -1018 -529 -994
rect -523 -1018 -495 -994
rect -589 -1110 -529 -1086
rect -523 -1110 -495 -1086
rect 151 -1128 211 -1104
rect 894 -1131 954 -1107
rect 1653 -1131 1713 -1107
rect 2389 -1131 2449 -1107
rect -159 -1176 -99 -1152
rect 78 -1176 138 -1152
rect -589 -1202 -529 -1178
rect -523 -1202 -495 -1178
rect 252 -1196 312 -1172
rect 584 -1179 644 -1155
rect 821 -1179 881 -1155
rect 995 -1199 1055 -1175
rect 1343 -1179 1403 -1155
rect 1580 -1179 1640 -1155
rect 1754 -1199 1814 -1175
rect 2079 -1179 2139 -1155
rect 2316 -1179 2376 -1155
rect 2490 -1199 2550 -1175
rect -232 -1224 -172 -1200
rect -58 -1244 2 -1220
rect 166 -1237 226 -1213
rect 511 -1227 571 -1203
rect 685 -1247 745 -1223
rect 909 -1240 969 -1216
rect 1270 -1227 1330 -1203
rect 1444 -1247 1504 -1223
rect 1668 -1240 1728 -1216
rect 2006 -1227 2066 -1203
rect 2180 -1247 2240 -1223
rect 2404 -1240 2464 -1216
rect -584 -1293 -524 -1269
rect -518 -1293 -490 -1269
rect -144 -1285 -84 -1261
rect 599 -1288 659 -1264
rect 1358 -1288 1418 -1264
rect 2094 -1288 2154 -1264
rect 138 -1343 198 -1319
rect 204 -1343 232 -1319
rect 297 -1343 357 -1319
rect 365 -1343 393 -1319
rect 881 -1346 941 -1322
rect 947 -1346 975 -1322
rect 1040 -1346 1100 -1322
rect 1108 -1346 1136 -1322
rect 1640 -1346 1700 -1322
rect 1706 -1346 1734 -1322
rect 1799 -1346 1859 -1322
rect 1867 -1346 1895 -1322
rect 2376 -1346 2436 -1322
rect 2442 -1346 2470 -1322
rect 2535 -1346 2595 -1322
rect 2603 -1346 2631 -1322
rect -587 -1385 -527 -1361
rect -521 -1385 -493 -1361
rect -173 -1394 -113 -1370
rect -107 -1394 -79 -1370
rect 570 -1397 630 -1373
rect 636 -1397 664 -1373
rect 1329 -1397 1389 -1373
rect 1395 -1397 1423 -1373
rect 2065 -1397 2125 -1373
rect 2131 -1397 2159 -1373
rect -587 -1477 -527 -1453
rect -521 -1477 -493 -1453
rect -587 -1569 -527 -1545
rect -521 -1569 -493 -1545
rect -586 -1689 -526 -1665
rect -520 -1689 -492 -1665
rect 7 -1745 67 -1721
rect 496 -1745 556 -1721
rect 880 -1745 940 -1721
rect -589 -1781 -529 -1757
rect -523 -1781 -495 -1757
rect 1295 -1769 1355 -1745
rect -66 -1793 -6 -1769
rect 108 -1813 168 -1789
rect 423 -1793 483 -1769
rect 234 -1817 262 -1793
rect 597 -1813 657 -1789
rect 807 -1793 867 -1769
rect 670 -1817 698 -1793
rect 1015 -1813 1075 -1789
rect 1088 -1817 1116 -1793
rect 1222 -1817 1282 -1793
rect -589 -1873 -529 -1849
rect -523 -1873 -495 -1849
rect 22 -1854 82 -1830
rect 511 -1854 571 -1830
rect 895 -1854 955 -1830
rect 1396 -1837 1456 -1813
rect 1464 -1837 1492 -1813
rect 1310 -1878 1370 -1854
rect -589 -1965 -529 -1941
rect -523 -1965 -495 -1941
rect -584 -2056 -524 -2032
rect -518 -2056 -486 -2032
rect 327 -2103 424 -2079
rect 435 -2103 463 -2079
rect 743 -2103 840 -2079
rect 851 -2103 879 -2079
rect 1193 -2103 1290 -2079
rect 1301 -2103 1329 -2079
rect -587 -2148 -527 -2124
rect -521 -2148 -493 -2124
rect 249 -2156 277 -2132
rect 665 -2156 693 -2132
rect 1109 -2156 1137 -2132
rect -40 -2180 -12 -2156
rect 47 -2188 107 -2164
rect 113 -2188 141 -2164
rect -587 -2240 -527 -2216
rect -521 -2240 -493 -2216
rect 249 -2248 277 -2224
rect 345 -2240 442 -2216
rect 453 -2240 481 -2216
rect -42 -2273 -14 -2249
rect 658 -2276 686 -2252
rect 761 -2268 858 -2244
rect 869 -2268 897 -2244
rect 1108 -2248 1136 -2224
rect 1211 -2240 1308 -2216
rect 1319 -2240 1347 -2216
rect 48 -2304 108 -2280
rect 114 -2304 142 -2280
rect 950 -2286 1010 -2262
rect 1016 -2286 1044 -2262
rect 1431 -2281 1547 -2257
rect 1555 -2281 1583 -2257
rect -587 -2332 -527 -2308
rect -521 -2332 -493 -2308
rect 541 -2325 601 -2301
rect 607 -2325 635 -2301
rect 29 -2482 152 -2458
rect 160 -2482 188 -2458
rect 299 -2482 422 -2458
rect 430 -2482 458 -2458
rect -586 -2616 -526 -2592
rect -520 -2616 -492 -2592
rect -589 -2708 -529 -2684
rect -523 -2708 -495 -2684
rect -88 -2775 -28 -2751
rect -22 -2775 6 -2751
rect -589 -2800 -529 -2776
rect -523 -2800 -495 -2776
rect -88 -2868 -28 -2844
rect -22 -2868 6 -2844
rect -589 -2892 -529 -2868
rect -523 -2892 -495 -2868
rect -584 -2983 -524 -2959
rect -518 -2983 -486 -2959
rect -88 -2960 -28 -2936
rect -22 -2960 6 -2936
rect -587 -3075 -527 -3051
rect -521 -3075 -493 -3051
rect -88 -3053 -28 -3029
rect -22 -3053 6 -3029
rect -587 -3167 -527 -3143
rect -521 -3167 -493 -3143
rect -587 -3259 -527 -3235
rect -521 -3259 -493 -3235
<< ntransistor >>
rect -872 100 -868 108
rect -796 94 -792 102
rect -775 94 -771 102
rect -730 94 -726 102
rect -626 94 -622 102
rect -605 94 -601 102
rect -560 94 -556 102
rect -869 -9 -865 -1
rect -796 -15 -792 -7
rect -775 -15 -771 -7
rect -730 -15 -726 -7
rect -630 -15 -626 -7
rect -609 -15 -605 -7
rect -564 -15 -560 -7
rect -436 -16 -432 -8
rect -147 -69 -143 -61
rect -126 -69 -122 -61
rect 451 -69 455 -61
rect 472 -69 476 -61
rect -220 -117 -216 -109
rect -199 -117 -195 -109
rect 1330 -69 1334 -61
rect 1351 -69 1355 -61
rect 378 -117 382 -109
rect 399 -117 403 -109
rect -574 -170 -570 -162
rect -553 -170 -549 -162
rect -508 -170 -504 -162
rect -46 -137 -42 -129
rect -25 -137 -21 -129
rect 2098 -69 2102 -61
rect 2119 -69 2123 -61
rect 1257 -117 1261 -109
rect 1278 -117 1282 -109
rect 552 -137 556 -129
rect 573 -137 577 -129
rect 2025 -117 2029 -109
rect 2046 -117 2050 -109
rect 1431 -137 1435 -129
rect 1452 -137 1456 -129
rect 2199 -137 2203 -129
rect 2220 -137 2224 -129
rect -132 -178 -128 -170
rect -111 -178 -107 -170
rect 466 -178 470 -170
rect 487 -178 491 -170
rect 1345 -178 1349 -170
rect 1366 -178 1370 -170
rect 2113 -178 2117 -170
rect 2134 -178 2138 -170
rect -577 -262 -573 -254
rect -556 -262 -552 -254
rect -511 -262 -507 -254
rect -577 -354 -573 -346
rect -556 -354 -552 -346
rect -511 -354 -507 -346
rect 134 -372 138 -364
rect 155 -372 159 -364
rect 877 -375 881 -367
rect 898 -375 902 -367
rect -176 -420 -172 -412
rect -155 -420 -151 -412
rect 61 -420 65 -412
rect 82 -420 86 -412
rect -577 -446 -573 -438
rect -556 -446 -552 -438
rect -511 -446 -507 -438
rect 1636 -375 1640 -367
rect 1657 -375 1661 -367
rect 567 -423 571 -415
rect 588 -423 592 -415
rect 804 -423 808 -415
rect 825 -423 829 -415
rect -249 -468 -245 -460
rect -228 -468 -224 -460
rect 235 -440 239 -432
rect 256 -440 260 -432
rect 2372 -375 2376 -367
rect 2393 -375 2397 -367
rect 1326 -423 1330 -415
rect 1347 -423 1351 -415
rect 1563 -423 1567 -415
rect 1584 -423 1588 -415
rect 494 -471 498 -463
rect 515 -471 519 -463
rect -75 -488 -71 -480
rect -54 -488 -50 -480
rect 149 -481 153 -473
rect 170 -481 174 -473
rect 978 -443 982 -435
rect 999 -443 1003 -435
rect 2062 -423 2066 -415
rect 2083 -423 2087 -415
rect 2299 -423 2303 -415
rect 2320 -423 2324 -415
rect 1253 -471 1257 -463
rect 1274 -471 1278 -463
rect -161 -529 -157 -521
rect -140 -529 -136 -521
rect 668 -491 672 -483
rect 689 -491 693 -483
rect 892 -484 896 -476
rect 913 -484 917 -476
rect 1737 -443 1741 -435
rect 1758 -443 1762 -435
rect 1989 -471 1993 -463
rect 2010 -471 2014 -463
rect 1427 -491 1431 -483
rect 1448 -491 1452 -483
rect 1651 -484 1655 -476
rect 1672 -484 1676 -476
rect 2473 -443 2477 -435
rect 2494 -443 2498 -435
rect 2163 -491 2167 -483
rect 2184 -491 2188 -483
rect 2387 -484 2391 -476
rect 2408 -484 2412 -476
rect -572 -537 -568 -529
rect -551 -537 -547 -529
rect -506 -537 -502 -529
rect 582 -532 586 -524
rect 603 -532 607 -524
rect 1341 -532 1345 -524
rect 1362 -532 1366 -524
rect 2077 -532 2081 -524
rect 2098 -532 2102 -524
rect 121 -587 125 -579
rect 142 -587 146 -579
rect 187 -587 191 -579
rect 280 -590 284 -582
rect 301 -590 305 -582
rect 348 -590 352 -582
rect -575 -629 -571 -621
rect -554 -629 -550 -621
rect -509 -629 -505 -621
rect 864 -590 868 -582
rect 885 -590 889 -582
rect 930 -590 934 -582
rect 1023 -593 1027 -585
rect 1044 -593 1048 -585
rect 1091 -593 1095 -585
rect 1623 -590 1627 -582
rect 1644 -590 1648 -582
rect 1689 -590 1693 -582
rect 1782 -593 1786 -585
rect 1803 -593 1807 -585
rect 1850 -593 1854 -585
rect 2359 -590 2363 -582
rect 2380 -590 2384 -582
rect 2425 -590 2429 -582
rect 2518 -593 2522 -585
rect 2539 -593 2543 -585
rect 2586 -593 2590 -585
rect -190 -638 -186 -630
rect -169 -638 -165 -630
rect -124 -638 -120 -630
rect 553 -641 557 -633
rect 574 -641 578 -633
rect 619 -641 623 -633
rect 1312 -641 1316 -633
rect 1333 -641 1337 -633
rect 1378 -641 1382 -633
rect 2048 -641 2052 -633
rect 2069 -641 2073 -633
rect 2114 -641 2118 -633
rect -575 -721 -571 -713
rect -554 -721 -550 -713
rect -509 -721 -505 -713
rect -575 -813 -571 -805
rect -554 -813 -550 -805
rect -509 -813 -505 -805
rect -118 -862 -114 -854
rect -97 -862 -93 -854
rect 480 -862 484 -854
rect 501 -862 505 -854
rect -191 -910 -187 -902
rect -170 -910 -166 -902
rect 1359 -862 1363 -854
rect 1380 -862 1384 -854
rect 407 -910 411 -902
rect 428 -910 432 -902
rect -574 -963 -570 -955
rect -553 -963 -549 -955
rect -508 -963 -504 -955
rect -17 -930 -13 -922
rect 4 -930 8 -922
rect 2127 -862 2131 -854
rect 2148 -862 2152 -854
rect 1286 -910 1290 -902
rect 1307 -910 1311 -902
rect 581 -930 585 -922
rect 602 -930 606 -922
rect 2054 -910 2058 -902
rect 2075 -910 2079 -902
rect 1460 -930 1464 -922
rect 1481 -930 1485 -922
rect 2228 -930 2232 -922
rect 2249 -930 2253 -922
rect -103 -971 -99 -963
rect -82 -971 -78 -963
rect 495 -971 499 -963
rect 516 -971 520 -963
rect 1374 -971 1378 -963
rect 1395 -971 1399 -963
rect 2142 -971 2146 -963
rect 2163 -971 2167 -963
rect -577 -1055 -573 -1047
rect -556 -1055 -552 -1047
rect -511 -1055 -507 -1047
rect -577 -1147 -573 -1139
rect -556 -1147 -552 -1139
rect -511 -1147 -507 -1139
rect 163 -1165 167 -1157
rect 184 -1165 188 -1157
rect 906 -1168 910 -1160
rect 927 -1168 931 -1160
rect -147 -1213 -143 -1205
rect -126 -1213 -122 -1205
rect 90 -1213 94 -1205
rect 111 -1213 115 -1205
rect -577 -1239 -573 -1231
rect -556 -1239 -552 -1231
rect -511 -1239 -507 -1231
rect 1665 -1168 1669 -1160
rect 1686 -1168 1690 -1160
rect 596 -1216 600 -1208
rect 617 -1216 621 -1208
rect 833 -1216 837 -1208
rect 854 -1216 858 -1208
rect -220 -1261 -216 -1253
rect -199 -1261 -195 -1253
rect 264 -1233 268 -1225
rect 285 -1233 289 -1225
rect 2401 -1168 2405 -1160
rect 2422 -1168 2426 -1160
rect 1355 -1216 1359 -1208
rect 1376 -1216 1380 -1208
rect 1592 -1216 1596 -1208
rect 1613 -1216 1617 -1208
rect 523 -1264 527 -1256
rect 544 -1264 548 -1256
rect -46 -1281 -42 -1273
rect -25 -1281 -21 -1273
rect 178 -1274 182 -1266
rect 199 -1274 203 -1266
rect 1007 -1236 1011 -1228
rect 1028 -1236 1032 -1228
rect 2091 -1216 2095 -1208
rect 2112 -1216 2116 -1208
rect 2328 -1216 2332 -1208
rect 2349 -1216 2353 -1208
rect 1282 -1264 1286 -1256
rect 1303 -1264 1307 -1256
rect -132 -1322 -128 -1314
rect -111 -1322 -107 -1314
rect 697 -1284 701 -1276
rect 718 -1284 722 -1276
rect 921 -1277 925 -1269
rect 942 -1277 946 -1269
rect 1766 -1236 1770 -1228
rect 1787 -1236 1791 -1228
rect 2018 -1264 2022 -1256
rect 2039 -1264 2043 -1256
rect 1456 -1284 1460 -1276
rect 1477 -1284 1481 -1276
rect 1680 -1277 1684 -1269
rect 1701 -1277 1705 -1269
rect 2502 -1236 2506 -1228
rect 2523 -1236 2527 -1228
rect 2192 -1284 2196 -1276
rect 2213 -1284 2217 -1276
rect 2416 -1277 2420 -1269
rect 2437 -1277 2441 -1269
rect -572 -1330 -568 -1322
rect -551 -1330 -547 -1322
rect -506 -1330 -502 -1322
rect 611 -1325 615 -1317
rect 632 -1325 636 -1317
rect 1370 -1325 1374 -1317
rect 1391 -1325 1395 -1317
rect 2106 -1325 2110 -1317
rect 2127 -1325 2131 -1317
rect 150 -1380 154 -1372
rect 171 -1380 175 -1372
rect 216 -1380 220 -1372
rect 309 -1383 313 -1375
rect 330 -1383 334 -1375
rect 377 -1383 381 -1375
rect -575 -1422 -571 -1414
rect -554 -1422 -550 -1414
rect -509 -1422 -505 -1414
rect 893 -1383 897 -1375
rect 914 -1383 918 -1375
rect 959 -1383 963 -1375
rect 1052 -1386 1056 -1378
rect 1073 -1386 1077 -1378
rect 1120 -1386 1124 -1378
rect 1652 -1383 1656 -1375
rect 1673 -1383 1677 -1375
rect 1718 -1383 1722 -1375
rect 1811 -1386 1815 -1378
rect 1832 -1386 1836 -1378
rect 1879 -1386 1883 -1378
rect 2388 -1383 2392 -1375
rect 2409 -1383 2413 -1375
rect 2454 -1383 2458 -1375
rect 2547 -1386 2551 -1378
rect 2568 -1386 2572 -1378
rect 2615 -1386 2619 -1378
rect -161 -1431 -157 -1423
rect -140 -1431 -136 -1423
rect -95 -1431 -91 -1423
rect 582 -1434 586 -1426
rect 603 -1434 607 -1426
rect 648 -1434 652 -1426
rect 1341 -1434 1345 -1426
rect 1362 -1434 1366 -1426
rect 1407 -1434 1411 -1426
rect 2077 -1434 2081 -1426
rect 2098 -1434 2102 -1426
rect 2143 -1434 2147 -1426
rect -575 -1514 -571 -1506
rect -554 -1514 -550 -1506
rect -509 -1514 -505 -1506
rect -575 -1606 -571 -1598
rect -554 -1606 -550 -1598
rect -509 -1606 -505 -1598
rect -574 -1726 -570 -1718
rect -553 -1726 -549 -1718
rect -508 -1726 -504 -1718
rect 19 -1782 23 -1774
rect 40 -1782 44 -1774
rect -577 -1818 -573 -1810
rect -556 -1818 -552 -1810
rect -511 -1818 -507 -1810
rect 508 -1782 512 -1774
rect 529 -1782 533 -1774
rect -54 -1830 -50 -1822
rect -33 -1830 -29 -1822
rect 892 -1782 896 -1774
rect 913 -1782 917 -1774
rect 435 -1830 439 -1822
rect 456 -1830 460 -1822
rect 120 -1850 124 -1842
rect 141 -1850 145 -1842
rect 246 -1848 250 -1840
rect 819 -1830 823 -1822
rect 840 -1830 844 -1822
rect 609 -1850 613 -1842
rect 630 -1850 634 -1842
rect 682 -1848 686 -1840
rect 1307 -1806 1311 -1798
rect 1328 -1806 1332 -1798
rect 1027 -1850 1031 -1842
rect 1048 -1850 1052 -1842
rect 1100 -1848 1104 -1840
rect 1234 -1854 1238 -1846
rect 1255 -1854 1259 -1846
rect 34 -1891 38 -1883
rect 55 -1891 59 -1883
rect 523 -1891 527 -1883
rect 544 -1891 548 -1883
rect 907 -1891 911 -1883
rect 928 -1891 932 -1883
rect -577 -1910 -573 -1902
rect -556 -1910 -552 -1902
rect -511 -1910 -507 -1902
rect 1408 -1874 1412 -1866
rect 1429 -1874 1433 -1866
rect 1476 -1868 1480 -1860
rect 1322 -1915 1326 -1907
rect 1343 -1915 1347 -1907
rect -577 -2002 -573 -1994
rect -556 -2002 -552 -1994
rect -511 -2002 -507 -1994
rect -572 -2093 -568 -2085
rect -551 -2093 -547 -2085
rect -506 -2093 -502 -2085
rect -575 -2185 -571 -2177
rect -554 -2185 -550 -2177
rect -509 -2185 -505 -2177
rect -28 -2211 -24 -2203
rect 339 -2169 343 -2161
rect 372 -2169 376 -2161
rect 396 -2169 400 -2161
rect 447 -2169 451 -2161
rect 755 -2169 759 -2161
rect 788 -2169 792 -2161
rect 812 -2169 816 -2161
rect 863 -2169 867 -2161
rect 1205 -2169 1209 -2161
rect 1238 -2169 1242 -2161
rect 1262 -2169 1266 -2161
rect 1313 -2169 1317 -2161
rect 261 -2193 265 -2185
rect 677 -2193 681 -2185
rect 1121 -2193 1125 -2185
rect 59 -2225 63 -2217
rect 80 -2225 84 -2217
rect 125 -2225 129 -2217
rect -575 -2277 -571 -2269
rect -554 -2277 -550 -2269
rect -509 -2277 -505 -2269
rect 261 -2285 265 -2277
rect -30 -2304 -26 -2296
rect 357 -2306 361 -2298
rect 390 -2306 394 -2298
rect 414 -2306 418 -2298
rect 465 -2306 469 -2298
rect 670 -2313 674 -2305
rect 60 -2341 64 -2333
rect 81 -2341 85 -2333
rect 126 -2341 130 -2333
rect 1120 -2285 1124 -2277
rect 1223 -2306 1227 -2298
rect 1256 -2306 1260 -2298
rect 1280 -2306 1284 -2298
rect 1331 -2306 1335 -2298
rect 962 -2323 966 -2315
rect 983 -2323 987 -2315
rect 1028 -2323 1032 -2315
rect 773 -2334 777 -2326
rect 806 -2334 810 -2326
rect 830 -2334 834 -2326
rect 881 -2334 885 -2326
rect 1443 -2335 1447 -2327
rect 1472 -2335 1476 -2327
rect 1496 -2335 1500 -2327
rect 1520 -2335 1524 -2327
rect 1567 -2335 1571 -2327
rect -575 -2369 -571 -2361
rect -554 -2369 -550 -2361
rect -509 -2369 -505 -2361
rect 553 -2362 557 -2354
rect 574 -2362 578 -2354
rect 619 -2362 623 -2354
rect 41 -2542 45 -2534
rect 62 -2542 66 -2534
rect 83 -2542 87 -2534
rect 104 -2542 108 -2534
rect 172 -2542 176 -2534
rect 311 -2545 315 -2537
rect 332 -2545 336 -2537
rect 353 -2545 357 -2537
rect 374 -2545 378 -2537
rect 442 -2545 446 -2537
rect -574 -2653 -570 -2645
rect -553 -2653 -549 -2645
rect -508 -2653 -504 -2645
rect -577 -2745 -573 -2737
rect -556 -2745 -552 -2737
rect -511 -2745 -507 -2737
rect -76 -2812 -72 -2804
rect -55 -2812 -51 -2804
rect -10 -2812 -6 -2804
rect -577 -2837 -573 -2829
rect -556 -2837 -552 -2829
rect -511 -2837 -507 -2829
rect -76 -2905 -72 -2897
rect -55 -2905 -51 -2897
rect -10 -2905 -6 -2897
rect -577 -2929 -573 -2921
rect -556 -2929 -552 -2921
rect -511 -2929 -507 -2921
rect -76 -2997 -72 -2989
rect -55 -2997 -51 -2989
rect -10 -2997 -6 -2989
rect -572 -3020 -568 -3012
rect -551 -3020 -547 -3012
rect -506 -3020 -502 -3012
rect -76 -3090 -72 -3082
rect -55 -3090 -51 -3082
rect -10 -3090 -6 -3082
rect -575 -3112 -571 -3104
rect -554 -3112 -550 -3104
rect -509 -3112 -505 -3104
rect -575 -3204 -571 -3196
rect -554 -3204 -550 -3196
rect -509 -3204 -505 -3196
rect -575 -3296 -571 -3288
rect -554 -3296 -550 -3288
rect -509 -3296 -505 -3288
<< ptransistor >>
rect -872 139 -868 147
rect -796 139 -792 147
rect -775 139 -771 147
rect -730 139 -726 147
rect -626 139 -622 147
rect -605 139 -601 147
rect -560 139 -556 147
rect -869 30 -865 38
rect -796 30 -792 38
rect -775 30 -771 38
rect -730 30 -726 38
rect -630 30 -626 38
rect -609 30 -605 38
rect -564 30 -560 38
rect -436 30 -432 38
rect -147 -24 -143 -16
rect -126 -24 -122 -16
rect 451 -24 455 -16
rect 472 -24 476 -16
rect 1330 -24 1334 -16
rect 1351 -24 1355 -16
rect 2098 -24 2102 -16
rect 2119 -24 2123 -16
rect -220 -72 -216 -64
rect -199 -72 -195 -64
rect 378 -72 382 -64
rect 399 -72 403 -64
rect -46 -92 -42 -84
rect -25 -92 -21 -84
rect -574 -125 -570 -117
rect -553 -125 -549 -117
rect -508 -125 -504 -117
rect -132 -133 -128 -125
rect -111 -133 -107 -125
rect 1257 -72 1261 -64
rect 1278 -72 1282 -64
rect 552 -92 556 -84
rect 573 -92 577 -84
rect 466 -133 470 -125
rect 487 -133 491 -125
rect 2025 -72 2029 -64
rect 2046 -72 2050 -64
rect 1431 -92 1435 -84
rect 1452 -92 1456 -84
rect 1345 -133 1349 -125
rect 1366 -133 1370 -125
rect 2199 -92 2203 -84
rect 2220 -92 2224 -84
rect 2113 -133 2117 -125
rect 2134 -133 2138 -125
rect -577 -217 -573 -209
rect -556 -217 -552 -209
rect -511 -217 -507 -209
rect -577 -309 -573 -301
rect -556 -309 -552 -301
rect -511 -309 -507 -301
rect 134 -327 138 -319
rect 155 -327 159 -319
rect 877 -330 881 -322
rect 898 -330 902 -322
rect 1636 -330 1640 -322
rect 1657 -330 1661 -322
rect 2372 -330 2376 -322
rect 2393 -330 2397 -322
rect -176 -375 -172 -367
rect -155 -375 -151 -367
rect 61 -375 65 -367
rect 82 -375 86 -367
rect -577 -401 -573 -393
rect -556 -401 -552 -393
rect -511 -401 -507 -393
rect 567 -378 571 -370
rect 588 -378 592 -370
rect 804 -378 808 -370
rect 825 -378 829 -370
rect 235 -395 239 -387
rect 256 -395 260 -387
rect -249 -423 -245 -415
rect -228 -423 -224 -415
rect -75 -443 -71 -435
rect -54 -443 -50 -435
rect 149 -436 153 -428
rect 170 -436 174 -428
rect 1326 -378 1330 -370
rect 1347 -378 1351 -370
rect 1563 -378 1567 -370
rect 1584 -378 1588 -370
rect 978 -398 982 -390
rect 999 -398 1003 -390
rect 494 -426 498 -418
rect 515 -426 519 -418
rect -161 -484 -157 -476
rect -140 -484 -136 -476
rect 668 -446 672 -438
rect 689 -446 693 -438
rect 892 -439 896 -431
rect 913 -439 917 -431
rect 2062 -378 2066 -370
rect 2083 -378 2087 -370
rect 2299 -378 2303 -370
rect 2320 -378 2324 -370
rect 1737 -398 1741 -390
rect 1758 -398 1762 -390
rect 1253 -426 1257 -418
rect 1274 -426 1278 -418
rect -572 -492 -568 -484
rect -551 -492 -547 -484
rect -506 -492 -502 -484
rect 582 -487 586 -479
rect 603 -487 607 -479
rect 1427 -446 1431 -438
rect 1448 -446 1452 -438
rect 1651 -439 1655 -431
rect 1672 -439 1676 -431
rect 2473 -398 2477 -390
rect 2494 -398 2498 -390
rect 1989 -426 1993 -418
rect 2010 -426 2014 -418
rect 1341 -487 1345 -479
rect 1362 -487 1366 -479
rect 2163 -446 2167 -438
rect 2184 -446 2188 -438
rect 2387 -439 2391 -431
rect 2408 -439 2412 -431
rect 2077 -487 2081 -479
rect 2098 -487 2102 -479
rect 121 -542 125 -534
rect 142 -542 146 -534
rect 187 -542 191 -534
rect 280 -542 284 -534
rect 301 -542 305 -534
rect 348 -542 352 -534
rect -575 -584 -571 -576
rect -554 -584 -550 -576
rect -509 -584 -505 -576
rect -190 -593 -186 -585
rect -169 -593 -165 -585
rect -124 -593 -120 -585
rect 864 -545 868 -537
rect 885 -545 889 -537
rect 930 -545 934 -537
rect 1023 -545 1027 -537
rect 1044 -545 1048 -537
rect 1091 -545 1095 -537
rect 1623 -545 1627 -537
rect 1644 -545 1648 -537
rect 1689 -545 1693 -537
rect 1782 -545 1786 -537
rect 1803 -545 1807 -537
rect 1850 -545 1854 -537
rect 2359 -545 2363 -537
rect 2380 -545 2384 -537
rect 2425 -545 2429 -537
rect 2518 -545 2522 -537
rect 2539 -545 2543 -537
rect 2586 -545 2590 -537
rect 553 -596 557 -588
rect 574 -596 578 -588
rect 619 -596 623 -588
rect 1312 -596 1316 -588
rect 1333 -596 1337 -588
rect 1378 -596 1382 -588
rect 2048 -596 2052 -588
rect 2069 -596 2073 -588
rect 2114 -596 2118 -588
rect -575 -676 -571 -668
rect -554 -676 -550 -668
rect -509 -676 -505 -668
rect -575 -768 -571 -760
rect -554 -768 -550 -760
rect -509 -768 -505 -760
rect -118 -817 -114 -809
rect -97 -817 -93 -809
rect 480 -817 484 -809
rect 501 -817 505 -809
rect 1359 -817 1363 -809
rect 1380 -817 1384 -809
rect 2127 -817 2131 -809
rect 2148 -817 2152 -809
rect -191 -865 -187 -857
rect -170 -865 -166 -857
rect 407 -865 411 -857
rect 428 -865 432 -857
rect -17 -885 -13 -877
rect 4 -885 8 -877
rect -574 -918 -570 -910
rect -553 -918 -549 -910
rect -508 -918 -504 -910
rect -103 -926 -99 -918
rect -82 -926 -78 -918
rect 1286 -865 1290 -857
rect 1307 -865 1311 -857
rect 581 -885 585 -877
rect 602 -885 606 -877
rect 495 -926 499 -918
rect 516 -926 520 -918
rect 2054 -865 2058 -857
rect 2075 -865 2079 -857
rect 1460 -885 1464 -877
rect 1481 -885 1485 -877
rect 1374 -926 1378 -918
rect 1395 -926 1399 -918
rect 2228 -885 2232 -877
rect 2249 -885 2253 -877
rect 2142 -926 2146 -918
rect 2163 -926 2167 -918
rect -577 -1010 -573 -1002
rect -556 -1010 -552 -1002
rect -511 -1010 -507 -1002
rect -577 -1102 -573 -1094
rect -556 -1102 -552 -1094
rect -511 -1102 -507 -1094
rect 163 -1120 167 -1112
rect 184 -1120 188 -1112
rect 906 -1123 910 -1115
rect 927 -1123 931 -1115
rect 1665 -1123 1669 -1115
rect 1686 -1123 1690 -1115
rect 2401 -1123 2405 -1115
rect 2422 -1123 2426 -1115
rect -147 -1168 -143 -1160
rect -126 -1168 -122 -1160
rect 90 -1168 94 -1160
rect 111 -1168 115 -1160
rect -577 -1194 -573 -1186
rect -556 -1194 -552 -1186
rect -511 -1194 -507 -1186
rect 596 -1171 600 -1163
rect 617 -1171 621 -1163
rect 833 -1171 837 -1163
rect 854 -1171 858 -1163
rect 264 -1188 268 -1180
rect 285 -1188 289 -1180
rect -220 -1216 -216 -1208
rect -199 -1216 -195 -1208
rect -46 -1236 -42 -1228
rect -25 -1236 -21 -1228
rect 178 -1229 182 -1221
rect 199 -1229 203 -1221
rect 1355 -1171 1359 -1163
rect 1376 -1171 1380 -1163
rect 1592 -1171 1596 -1163
rect 1613 -1171 1617 -1163
rect 1007 -1191 1011 -1183
rect 1028 -1191 1032 -1183
rect 523 -1219 527 -1211
rect 544 -1219 548 -1211
rect -132 -1277 -128 -1269
rect -111 -1277 -107 -1269
rect 697 -1239 701 -1231
rect 718 -1239 722 -1231
rect 921 -1232 925 -1224
rect 942 -1232 946 -1224
rect 2091 -1171 2095 -1163
rect 2112 -1171 2116 -1163
rect 2328 -1171 2332 -1163
rect 2349 -1171 2353 -1163
rect 1766 -1191 1770 -1183
rect 1787 -1191 1791 -1183
rect 1282 -1219 1286 -1211
rect 1303 -1219 1307 -1211
rect -572 -1285 -568 -1277
rect -551 -1285 -547 -1277
rect -506 -1285 -502 -1277
rect 611 -1280 615 -1272
rect 632 -1280 636 -1272
rect 1456 -1239 1460 -1231
rect 1477 -1239 1481 -1231
rect 1680 -1232 1684 -1224
rect 1701 -1232 1705 -1224
rect 2502 -1191 2506 -1183
rect 2523 -1191 2527 -1183
rect 2018 -1219 2022 -1211
rect 2039 -1219 2043 -1211
rect 1370 -1280 1374 -1272
rect 1391 -1280 1395 -1272
rect 2192 -1239 2196 -1231
rect 2213 -1239 2217 -1231
rect 2416 -1232 2420 -1224
rect 2437 -1232 2441 -1224
rect 2106 -1280 2110 -1272
rect 2127 -1280 2131 -1272
rect 150 -1335 154 -1327
rect 171 -1335 175 -1327
rect 216 -1335 220 -1327
rect 309 -1335 313 -1327
rect 330 -1335 334 -1327
rect 377 -1335 381 -1327
rect -575 -1377 -571 -1369
rect -554 -1377 -550 -1369
rect -509 -1377 -505 -1369
rect -161 -1386 -157 -1378
rect -140 -1386 -136 -1378
rect -95 -1386 -91 -1378
rect 893 -1338 897 -1330
rect 914 -1338 918 -1330
rect 959 -1338 963 -1330
rect 1052 -1338 1056 -1330
rect 1073 -1338 1077 -1330
rect 1120 -1338 1124 -1330
rect 1652 -1338 1656 -1330
rect 1673 -1338 1677 -1330
rect 1718 -1338 1722 -1330
rect 1811 -1338 1815 -1330
rect 1832 -1338 1836 -1330
rect 1879 -1338 1883 -1330
rect 2388 -1338 2392 -1330
rect 2409 -1338 2413 -1330
rect 2454 -1338 2458 -1330
rect 2547 -1338 2551 -1330
rect 2568 -1338 2572 -1330
rect 2615 -1338 2619 -1330
rect 582 -1389 586 -1381
rect 603 -1389 607 -1381
rect 648 -1389 652 -1381
rect 1341 -1389 1345 -1381
rect 1362 -1389 1366 -1381
rect 1407 -1389 1411 -1381
rect 2077 -1389 2081 -1381
rect 2098 -1389 2102 -1381
rect 2143 -1389 2147 -1381
rect -575 -1469 -571 -1461
rect -554 -1469 -550 -1461
rect -509 -1469 -505 -1461
rect -575 -1561 -571 -1553
rect -554 -1561 -550 -1553
rect -509 -1561 -505 -1553
rect -574 -1681 -570 -1673
rect -553 -1681 -549 -1673
rect -508 -1681 -504 -1673
rect 19 -1737 23 -1729
rect 40 -1737 44 -1729
rect 508 -1737 512 -1729
rect 529 -1737 533 -1729
rect 892 -1737 896 -1729
rect 913 -1737 917 -1729
rect -577 -1773 -573 -1765
rect -556 -1773 -552 -1765
rect -511 -1773 -507 -1765
rect 1307 -1761 1311 -1753
rect 1328 -1761 1332 -1753
rect -54 -1785 -50 -1777
rect -33 -1785 -29 -1777
rect 435 -1785 439 -1777
rect 456 -1785 460 -1777
rect 120 -1805 124 -1797
rect 141 -1805 145 -1797
rect 34 -1846 38 -1838
rect 55 -1846 59 -1838
rect 246 -1809 250 -1801
rect 819 -1785 823 -1777
rect 840 -1785 844 -1777
rect 609 -1805 613 -1797
rect 630 -1805 634 -1797
rect -577 -1865 -573 -1857
rect -556 -1865 -552 -1857
rect -511 -1865 -507 -1857
rect 523 -1846 527 -1838
rect 544 -1846 548 -1838
rect 682 -1809 686 -1801
rect 1027 -1805 1031 -1797
rect 1048 -1805 1052 -1797
rect 907 -1846 911 -1838
rect 928 -1846 932 -1838
rect 1100 -1809 1104 -1801
rect 1234 -1809 1238 -1801
rect 1255 -1809 1259 -1801
rect 1408 -1829 1412 -1821
rect 1429 -1829 1433 -1821
rect 1476 -1829 1480 -1821
rect 1322 -1870 1326 -1862
rect 1343 -1870 1347 -1862
rect -577 -1957 -573 -1949
rect -556 -1957 -552 -1949
rect -511 -1957 -507 -1949
rect -572 -2048 -568 -2040
rect -551 -2048 -547 -2040
rect -506 -2048 -502 -2040
rect 339 -2095 343 -2087
rect 372 -2095 376 -2087
rect 396 -2095 400 -2087
rect 447 -2095 451 -2087
rect 755 -2095 759 -2087
rect 788 -2095 792 -2087
rect 812 -2095 816 -2087
rect 863 -2095 867 -2087
rect 1205 -2095 1209 -2087
rect 1238 -2095 1242 -2087
rect 1262 -2095 1266 -2087
rect 1313 -2095 1317 -2087
rect -575 -2140 -571 -2132
rect -554 -2140 -550 -2132
rect -509 -2140 -505 -2132
rect 261 -2148 265 -2140
rect -28 -2172 -24 -2164
rect 59 -2180 63 -2172
rect 80 -2180 84 -2172
rect 125 -2180 129 -2172
rect 677 -2148 681 -2140
rect 1121 -2148 1125 -2140
rect -575 -2232 -571 -2224
rect -554 -2232 -550 -2224
rect -509 -2232 -505 -2224
rect 357 -2232 361 -2224
rect 390 -2232 394 -2224
rect 414 -2232 418 -2224
rect 465 -2232 469 -2224
rect 261 -2240 265 -2232
rect -30 -2265 -26 -2257
rect 60 -2296 64 -2288
rect 81 -2296 85 -2288
rect 126 -2296 130 -2288
rect -575 -2324 -571 -2316
rect -554 -2324 -550 -2316
rect -509 -2324 -505 -2316
rect 1223 -2232 1227 -2224
rect 1256 -2232 1260 -2224
rect 1280 -2232 1284 -2224
rect 1331 -2232 1335 -2224
rect 1120 -2240 1124 -2232
rect 773 -2260 777 -2252
rect 806 -2260 810 -2252
rect 830 -2260 834 -2252
rect 881 -2260 885 -2252
rect 670 -2268 674 -2260
rect 553 -2317 557 -2309
rect 574 -2317 578 -2309
rect 619 -2317 623 -2309
rect 962 -2278 966 -2270
rect 983 -2278 987 -2270
rect 1028 -2278 1032 -2270
rect 1443 -2273 1447 -2265
rect 1472 -2273 1476 -2265
rect 1496 -2273 1500 -2265
rect 1520 -2273 1524 -2265
rect 1567 -2273 1571 -2265
rect 41 -2474 45 -2466
rect 62 -2474 66 -2466
rect 83 -2474 87 -2466
rect 104 -2474 108 -2466
rect 172 -2474 176 -2466
rect 311 -2474 315 -2466
rect 332 -2474 336 -2466
rect 353 -2474 357 -2466
rect 374 -2474 378 -2466
rect 442 -2474 446 -2466
rect -574 -2608 -570 -2600
rect -553 -2608 -549 -2600
rect -508 -2608 -504 -2600
rect -577 -2700 -573 -2692
rect -556 -2700 -552 -2692
rect -511 -2700 -507 -2692
rect -76 -2767 -72 -2759
rect -55 -2767 -51 -2759
rect -10 -2767 -6 -2759
rect -577 -2792 -573 -2784
rect -556 -2792 -552 -2784
rect -511 -2792 -507 -2784
rect -76 -2860 -72 -2852
rect -55 -2860 -51 -2852
rect -10 -2860 -6 -2852
rect -577 -2884 -573 -2876
rect -556 -2884 -552 -2876
rect -511 -2884 -507 -2876
rect -76 -2952 -72 -2944
rect -55 -2952 -51 -2944
rect -10 -2952 -6 -2944
rect -572 -2975 -568 -2967
rect -551 -2975 -547 -2967
rect -506 -2975 -502 -2967
rect -76 -3045 -72 -3037
rect -55 -3045 -51 -3037
rect -10 -3045 -6 -3037
rect -575 -3067 -571 -3059
rect -554 -3067 -550 -3059
rect -509 -3067 -505 -3059
rect -575 -3159 -571 -3151
rect -554 -3159 -550 -3151
rect -509 -3159 -505 -3151
rect -575 -3251 -571 -3243
rect -554 -3251 -550 -3243
rect -509 -3251 -505 -3243
<< ndiffusion >>
rect -878 106 -872 108
rect -878 102 -877 106
rect -873 102 -872 106
rect -878 100 -872 102
rect -868 106 -862 108
rect -868 102 -867 106
rect -863 102 -862 106
rect -868 100 -862 102
rect -802 100 -796 102
rect -802 96 -801 100
rect -797 96 -796 100
rect -802 94 -796 96
rect -792 94 -775 102
rect -771 100 -754 102
rect -771 96 -768 100
rect -764 96 -754 100
rect -771 94 -754 96
rect -736 100 -730 102
rect -736 96 -735 100
rect -731 96 -730 100
rect -736 94 -730 96
rect -726 100 -720 102
rect -726 96 -725 100
rect -721 96 -720 100
rect -726 94 -720 96
rect -632 100 -626 102
rect -632 96 -631 100
rect -627 96 -626 100
rect -632 94 -626 96
rect -622 94 -605 102
rect -601 100 -584 102
rect -601 96 -598 100
rect -594 96 -584 100
rect -601 94 -584 96
rect -566 100 -560 102
rect -566 96 -565 100
rect -561 96 -560 100
rect -566 94 -560 96
rect -556 100 -550 102
rect -556 96 -555 100
rect -551 96 -550 100
rect -556 94 -550 96
rect -875 -3 -869 -1
rect -875 -7 -874 -3
rect -870 -7 -869 -3
rect -875 -9 -869 -7
rect -865 -3 -859 -1
rect -865 -7 -864 -3
rect -860 -7 -859 -3
rect -865 -9 -859 -7
rect -802 -9 -796 -7
rect -802 -13 -801 -9
rect -797 -13 -796 -9
rect -802 -15 -796 -13
rect -792 -15 -775 -7
rect -771 -9 -754 -7
rect -771 -13 -768 -9
rect -764 -13 -754 -9
rect -771 -15 -754 -13
rect -736 -9 -730 -7
rect -736 -13 -735 -9
rect -731 -13 -730 -9
rect -736 -15 -730 -13
rect -726 -9 -720 -7
rect -726 -13 -725 -9
rect -721 -13 -720 -9
rect -726 -15 -720 -13
rect -636 -9 -630 -7
rect -636 -13 -635 -9
rect -631 -13 -630 -9
rect -636 -15 -630 -13
rect -626 -15 -609 -7
rect -605 -9 -588 -7
rect -605 -13 -602 -9
rect -598 -13 -588 -9
rect -605 -15 -588 -13
rect -570 -9 -564 -7
rect -570 -13 -569 -9
rect -565 -13 -564 -9
rect -570 -15 -564 -13
rect -560 -9 -554 -7
rect -560 -13 -559 -9
rect -555 -13 -554 -9
rect -560 -15 -554 -13
rect -442 -10 -436 -8
rect -442 -14 -441 -10
rect -437 -14 -436 -10
rect -442 -16 -436 -14
rect -432 -10 -426 -8
rect -432 -14 -431 -10
rect -427 -14 -426 -10
rect -432 -16 -426 -14
rect -153 -63 -147 -61
rect -153 -67 -152 -63
rect -148 -67 -147 -63
rect -153 -69 -147 -67
rect -143 -69 -126 -61
rect -122 -63 -105 -61
rect -122 -67 -119 -63
rect -115 -67 -105 -63
rect 445 -63 451 -61
rect -122 -69 -105 -67
rect 445 -67 446 -63
rect 450 -67 451 -63
rect 445 -69 451 -67
rect 455 -69 472 -61
rect 476 -63 493 -61
rect 476 -67 479 -63
rect 483 -67 493 -63
rect 1324 -63 1330 -61
rect 476 -69 493 -67
rect -226 -111 -220 -109
rect -226 -115 -225 -111
rect -221 -115 -220 -111
rect -226 -117 -220 -115
rect -216 -117 -199 -109
rect -195 -111 -178 -109
rect -195 -115 -192 -111
rect -188 -115 -178 -111
rect -195 -117 -178 -115
rect 1324 -67 1325 -63
rect 1329 -67 1330 -63
rect 1324 -69 1330 -67
rect 1334 -69 1351 -61
rect 1355 -63 1372 -61
rect 1355 -67 1358 -63
rect 1362 -67 1372 -63
rect 2092 -63 2098 -61
rect 1355 -69 1372 -67
rect 372 -111 378 -109
rect 372 -115 373 -111
rect 377 -115 378 -111
rect 372 -117 378 -115
rect 382 -117 399 -109
rect 403 -111 420 -109
rect 403 -115 406 -111
rect 410 -115 420 -111
rect 403 -117 420 -115
rect -52 -131 -46 -129
rect -580 -164 -574 -162
rect -580 -168 -579 -164
rect -575 -168 -574 -164
rect -580 -170 -574 -168
rect -570 -170 -553 -162
rect -549 -164 -532 -162
rect -549 -168 -546 -164
rect -542 -168 -532 -164
rect -549 -170 -532 -168
rect -514 -164 -508 -162
rect -514 -168 -513 -164
rect -509 -168 -508 -164
rect -514 -170 -508 -168
rect -504 -164 -498 -162
rect -504 -168 -503 -164
rect -499 -168 -498 -164
rect -504 -170 -498 -168
rect -52 -135 -51 -131
rect -47 -135 -46 -131
rect -52 -137 -46 -135
rect -42 -137 -25 -129
rect -21 -131 -4 -129
rect -21 -135 -18 -131
rect -14 -135 -4 -131
rect 2092 -67 2093 -63
rect 2097 -67 2098 -63
rect 2092 -69 2098 -67
rect 2102 -69 2119 -61
rect 2123 -63 2140 -61
rect 2123 -67 2126 -63
rect 2130 -67 2140 -63
rect 2123 -69 2140 -67
rect 1251 -111 1257 -109
rect 1251 -115 1252 -111
rect 1256 -115 1257 -111
rect 1251 -117 1257 -115
rect 1261 -117 1278 -109
rect 1282 -111 1299 -109
rect 1282 -115 1285 -111
rect 1289 -115 1299 -111
rect 1282 -117 1299 -115
rect 546 -131 552 -129
rect -21 -137 -4 -135
rect 546 -135 547 -131
rect 551 -135 552 -131
rect 546 -137 552 -135
rect 556 -137 573 -129
rect 577 -131 594 -129
rect 577 -135 580 -131
rect 584 -135 594 -131
rect 2019 -111 2025 -109
rect 2019 -115 2020 -111
rect 2024 -115 2025 -111
rect 2019 -117 2025 -115
rect 2029 -117 2046 -109
rect 2050 -111 2067 -109
rect 2050 -115 2053 -111
rect 2057 -115 2067 -111
rect 2050 -117 2067 -115
rect 1425 -131 1431 -129
rect 577 -137 594 -135
rect 1425 -135 1426 -131
rect 1430 -135 1431 -131
rect 1425 -137 1431 -135
rect 1435 -137 1452 -129
rect 1456 -131 1473 -129
rect 1456 -135 1459 -131
rect 1463 -135 1473 -131
rect 2193 -131 2199 -129
rect 1456 -137 1473 -135
rect 2193 -135 2194 -131
rect 2198 -135 2199 -131
rect 2193 -137 2199 -135
rect 2203 -137 2220 -129
rect 2224 -131 2241 -129
rect 2224 -135 2227 -131
rect 2231 -135 2241 -131
rect 2224 -137 2241 -135
rect -138 -172 -132 -170
rect -138 -176 -137 -172
rect -133 -176 -132 -172
rect -138 -178 -132 -176
rect -128 -178 -111 -170
rect -107 -172 -90 -170
rect -107 -176 -104 -172
rect -100 -176 -90 -172
rect -107 -178 -90 -176
rect 460 -172 466 -170
rect 460 -176 461 -172
rect 465 -176 466 -172
rect 460 -178 466 -176
rect 470 -178 487 -170
rect 491 -172 508 -170
rect 491 -176 494 -172
rect 498 -176 508 -172
rect 491 -178 508 -176
rect 1339 -172 1345 -170
rect 1339 -176 1340 -172
rect 1344 -176 1345 -172
rect 1339 -178 1345 -176
rect 1349 -178 1366 -170
rect 1370 -172 1387 -170
rect 1370 -176 1373 -172
rect 1377 -176 1387 -172
rect 1370 -178 1387 -176
rect 2107 -172 2113 -170
rect 2107 -176 2108 -172
rect 2112 -176 2113 -172
rect 2107 -178 2113 -176
rect 2117 -178 2134 -170
rect 2138 -172 2155 -170
rect 2138 -176 2141 -172
rect 2145 -176 2155 -172
rect 2138 -178 2155 -176
rect -583 -256 -577 -254
rect -583 -260 -582 -256
rect -578 -260 -577 -256
rect -583 -262 -577 -260
rect -573 -262 -556 -254
rect -552 -256 -535 -254
rect -552 -260 -549 -256
rect -545 -260 -535 -256
rect -552 -262 -535 -260
rect -517 -256 -511 -254
rect -517 -260 -516 -256
rect -512 -260 -511 -256
rect -517 -262 -511 -260
rect -507 -256 -501 -254
rect -507 -260 -506 -256
rect -502 -260 -501 -256
rect -507 -262 -501 -260
rect -583 -348 -577 -346
rect -583 -352 -582 -348
rect -578 -352 -577 -348
rect -583 -354 -577 -352
rect -573 -354 -556 -346
rect -552 -348 -535 -346
rect -552 -352 -549 -348
rect -545 -352 -535 -348
rect -552 -354 -535 -352
rect -517 -348 -511 -346
rect -517 -352 -516 -348
rect -512 -352 -511 -348
rect -517 -354 -511 -352
rect -507 -348 -501 -346
rect -507 -352 -506 -348
rect -502 -352 -501 -348
rect -507 -354 -501 -352
rect 128 -366 134 -364
rect 128 -370 129 -366
rect 133 -370 134 -366
rect 128 -372 134 -370
rect 138 -372 155 -364
rect 159 -366 176 -364
rect 159 -370 162 -366
rect 166 -370 176 -366
rect 871 -369 877 -367
rect 159 -372 176 -370
rect 871 -373 872 -369
rect 876 -373 877 -369
rect 871 -375 877 -373
rect 881 -375 898 -367
rect 902 -369 919 -367
rect 902 -373 905 -369
rect 909 -373 919 -369
rect 1630 -369 1636 -367
rect 902 -375 919 -373
rect -182 -414 -176 -412
rect -182 -418 -181 -414
rect -177 -418 -176 -414
rect -182 -420 -176 -418
rect -172 -420 -155 -412
rect -151 -414 -134 -412
rect -151 -418 -148 -414
rect -144 -418 -134 -414
rect -151 -420 -134 -418
rect 55 -414 61 -412
rect 55 -418 56 -414
rect 60 -418 61 -414
rect 55 -420 61 -418
rect 65 -420 82 -412
rect 86 -414 103 -412
rect 86 -418 89 -414
rect 93 -418 103 -414
rect 86 -420 103 -418
rect -583 -440 -577 -438
rect -583 -444 -582 -440
rect -578 -444 -577 -440
rect -583 -446 -577 -444
rect -573 -446 -556 -438
rect -552 -440 -535 -438
rect -552 -444 -549 -440
rect -545 -444 -535 -440
rect -552 -446 -535 -444
rect -517 -440 -511 -438
rect -517 -444 -516 -440
rect -512 -444 -511 -440
rect -517 -446 -511 -444
rect -507 -440 -501 -438
rect -507 -444 -506 -440
rect -502 -444 -501 -440
rect -507 -446 -501 -444
rect 1630 -373 1631 -369
rect 1635 -373 1636 -369
rect 1630 -375 1636 -373
rect 1640 -375 1657 -367
rect 1661 -369 1678 -367
rect 1661 -373 1664 -369
rect 1668 -373 1678 -369
rect 2366 -369 2372 -367
rect 1661 -375 1678 -373
rect 561 -417 567 -415
rect 561 -421 562 -417
rect 566 -421 567 -417
rect 561 -423 567 -421
rect 571 -423 588 -415
rect 592 -417 609 -415
rect 592 -421 595 -417
rect 599 -421 609 -417
rect 592 -423 609 -421
rect 798 -417 804 -415
rect 798 -421 799 -417
rect 803 -421 804 -417
rect 798 -423 804 -421
rect 808 -423 825 -415
rect 829 -417 846 -415
rect 829 -421 832 -417
rect 836 -421 846 -417
rect 829 -423 846 -421
rect 229 -434 235 -432
rect -255 -462 -249 -460
rect -255 -466 -254 -462
rect -250 -466 -249 -462
rect -255 -468 -249 -466
rect -245 -468 -228 -460
rect -224 -462 -207 -460
rect -224 -466 -221 -462
rect -217 -466 -207 -462
rect -224 -468 -207 -466
rect 229 -438 230 -434
rect 234 -438 235 -434
rect 229 -440 235 -438
rect 239 -440 256 -432
rect 260 -434 277 -432
rect 260 -438 263 -434
rect 267 -438 277 -434
rect 260 -440 277 -438
rect 2366 -373 2367 -369
rect 2371 -373 2372 -369
rect 2366 -375 2372 -373
rect 2376 -375 2393 -367
rect 2397 -369 2414 -367
rect 2397 -373 2400 -369
rect 2404 -373 2414 -369
rect 2397 -375 2414 -373
rect 1320 -417 1326 -415
rect 1320 -421 1321 -417
rect 1325 -421 1326 -417
rect 1320 -423 1326 -421
rect 1330 -423 1347 -415
rect 1351 -417 1368 -415
rect 1351 -421 1354 -417
rect 1358 -421 1368 -417
rect 1351 -423 1368 -421
rect 1557 -417 1563 -415
rect 1557 -421 1558 -417
rect 1562 -421 1563 -417
rect 1557 -423 1563 -421
rect 1567 -423 1584 -415
rect 1588 -417 1605 -415
rect 1588 -421 1591 -417
rect 1595 -421 1605 -417
rect 1588 -423 1605 -421
rect 972 -437 978 -435
rect 488 -465 494 -463
rect 488 -469 489 -465
rect 493 -469 494 -465
rect 488 -471 494 -469
rect 498 -471 515 -463
rect 519 -465 536 -463
rect 519 -469 522 -465
rect 526 -469 536 -465
rect 519 -471 536 -469
rect 143 -475 149 -473
rect 143 -479 144 -475
rect 148 -479 149 -475
rect -81 -482 -75 -480
rect -81 -486 -80 -482
rect -76 -486 -75 -482
rect -81 -488 -75 -486
rect -71 -488 -54 -480
rect -50 -482 -33 -480
rect 143 -481 149 -479
rect 153 -481 170 -473
rect 174 -475 191 -473
rect 174 -479 177 -475
rect 181 -479 191 -475
rect 174 -481 191 -479
rect -50 -486 -47 -482
rect -43 -486 -33 -482
rect -50 -488 -33 -486
rect 972 -441 973 -437
rect 977 -441 978 -437
rect 972 -443 978 -441
rect 982 -443 999 -435
rect 1003 -437 1020 -435
rect 1003 -441 1006 -437
rect 1010 -441 1020 -437
rect 1003 -443 1020 -441
rect 2056 -417 2062 -415
rect 2056 -421 2057 -417
rect 2061 -421 2062 -417
rect 2056 -423 2062 -421
rect 2066 -423 2083 -415
rect 2087 -417 2104 -415
rect 2087 -421 2090 -417
rect 2094 -421 2104 -417
rect 2087 -423 2104 -421
rect 2293 -417 2299 -415
rect 2293 -421 2294 -417
rect 2298 -421 2299 -417
rect 2293 -423 2299 -421
rect 2303 -423 2320 -415
rect 2324 -417 2341 -415
rect 2324 -421 2327 -417
rect 2331 -421 2341 -417
rect 2324 -423 2341 -421
rect 1731 -437 1737 -435
rect 1247 -465 1253 -463
rect 1247 -469 1248 -465
rect 1252 -469 1253 -465
rect 1247 -471 1253 -469
rect 1257 -471 1274 -463
rect 1278 -465 1295 -463
rect 1278 -469 1281 -465
rect 1285 -469 1295 -465
rect 1278 -471 1295 -469
rect 886 -478 892 -476
rect 886 -482 887 -478
rect 891 -482 892 -478
rect 662 -485 668 -483
rect -167 -523 -161 -521
rect -167 -527 -166 -523
rect -162 -527 -161 -523
rect -167 -529 -161 -527
rect -157 -529 -140 -521
rect -136 -523 -119 -521
rect -136 -527 -133 -523
rect -129 -527 -119 -523
rect 662 -489 663 -485
rect 667 -489 668 -485
rect 662 -491 668 -489
rect 672 -491 689 -483
rect 693 -485 710 -483
rect 886 -484 892 -482
rect 896 -484 913 -476
rect 917 -478 934 -476
rect 917 -482 920 -478
rect 924 -482 934 -478
rect 917 -484 934 -482
rect 693 -489 696 -485
rect 700 -489 710 -485
rect 693 -491 710 -489
rect 1731 -441 1732 -437
rect 1736 -441 1737 -437
rect 1731 -443 1737 -441
rect 1741 -443 1758 -435
rect 1762 -437 1779 -435
rect 1762 -441 1765 -437
rect 1769 -441 1779 -437
rect 1762 -443 1779 -441
rect 2467 -437 2473 -435
rect 1983 -465 1989 -463
rect 1983 -469 1984 -465
rect 1988 -469 1989 -465
rect 1983 -471 1989 -469
rect 1993 -471 2010 -463
rect 2014 -465 2031 -463
rect 2014 -469 2017 -465
rect 2021 -469 2031 -465
rect 2014 -471 2031 -469
rect 1645 -478 1651 -476
rect 1645 -482 1646 -478
rect 1650 -482 1651 -478
rect 1421 -485 1427 -483
rect 1421 -489 1422 -485
rect 1426 -489 1427 -485
rect 1421 -491 1427 -489
rect 1431 -491 1448 -483
rect 1452 -485 1469 -483
rect 1645 -484 1651 -482
rect 1655 -484 1672 -476
rect 1676 -478 1693 -476
rect 1676 -482 1679 -478
rect 1683 -482 1693 -478
rect 1676 -484 1693 -482
rect 1452 -489 1455 -485
rect 1459 -489 1469 -485
rect 1452 -491 1469 -489
rect 2467 -441 2468 -437
rect 2472 -441 2473 -437
rect 2467 -443 2473 -441
rect 2477 -443 2494 -435
rect 2498 -437 2515 -435
rect 2498 -441 2501 -437
rect 2505 -441 2515 -437
rect 2498 -443 2515 -441
rect 2381 -478 2387 -476
rect 2381 -482 2382 -478
rect 2386 -482 2387 -478
rect 2157 -485 2163 -483
rect 2157 -489 2158 -485
rect 2162 -489 2163 -485
rect 2157 -491 2163 -489
rect 2167 -491 2184 -483
rect 2188 -485 2205 -483
rect 2381 -484 2387 -482
rect 2391 -484 2408 -476
rect 2412 -478 2429 -476
rect 2412 -482 2415 -478
rect 2419 -482 2429 -478
rect 2412 -484 2429 -482
rect 2188 -489 2191 -485
rect 2195 -489 2205 -485
rect 2188 -491 2205 -489
rect -136 -529 -119 -527
rect 576 -526 582 -524
rect -578 -531 -572 -529
rect -578 -535 -577 -531
rect -573 -535 -572 -531
rect -578 -537 -572 -535
rect -568 -537 -551 -529
rect -547 -531 -530 -529
rect -547 -535 -544 -531
rect -540 -535 -530 -531
rect -547 -537 -530 -535
rect -512 -531 -506 -529
rect -512 -535 -511 -531
rect -507 -535 -506 -531
rect -512 -537 -506 -535
rect -502 -531 -496 -529
rect -502 -535 -501 -531
rect -497 -535 -496 -531
rect -502 -537 -496 -535
rect 576 -530 577 -526
rect 581 -530 582 -526
rect 576 -532 582 -530
rect 586 -532 603 -524
rect 607 -526 624 -524
rect 607 -530 610 -526
rect 614 -530 624 -526
rect 607 -532 624 -530
rect 1335 -526 1341 -524
rect 1335 -530 1336 -526
rect 1340 -530 1341 -526
rect 1335 -532 1341 -530
rect 1345 -532 1362 -524
rect 1366 -526 1383 -524
rect 1366 -530 1369 -526
rect 1373 -530 1383 -526
rect 1366 -532 1383 -530
rect 2071 -526 2077 -524
rect 2071 -530 2072 -526
rect 2076 -530 2077 -526
rect 2071 -532 2077 -530
rect 2081 -532 2098 -524
rect 2102 -526 2119 -524
rect 2102 -530 2105 -526
rect 2109 -530 2119 -526
rect 2102 -532 2119 -530
rect 115 -581 121 -579
rect 115 -585 116 -581
rect 120 -585 121 -581
rect 115 -587 121 -585
rect 125 -587 142 -579
rect 146 -581 163 -579
rect 146 -585 149 -581
rect 153 -585 163 -581
rect 146 -587 163 -585
rect 181 -581 187 -579
rect 181 -585 182 -581
rect 186 -585 187 -581
rect 181 -587 187 -585
rect 191 -581 197 -579
rect 191 -585 192 -581
rect 196 -585 197 -581
rect 191 -587 197 -585
rect 274 -584 280 -582
rect 274 -588 275 -584
rect 279 -588 280 -584
rect 274 -590 280 -588
rect 284 -584 301 -582
rect 284 -588 285 -584
rect 289 -588 301 -584
rect 284 -590 301 -588
rect 305 -584 322 -582
rect 305 -588 308 -584
rect 312 -588 322 -584
rect 305 -590 322 -588
rect 342 -584 348 -582
rect 342 -588 343 -584
rect 347 -588 348 -584
rect 342 -590 348 -588
rect 352 -584 358 -582
rect 352 -588 353 -584
rect 357 -588 358 -584
rect 858 -584 864 -582
rect 858 -588 859 -584
rect 863 -588 864 -584
rect 352 -590 358 -588
rect -581 -623 -575 -621
rect -581 -627 -580 -623
rect -576 -627 -575 -623
rect -581 -629 -575 -627
rect -571 -629 -554 -621
rect -550 -623 -533 -621
rect -550 -627 -547 -623
rect -543 -627 -533 -623
rect -550 -629 -533 -627
rect -515 -623 -509 -621
rect -515 -627 -514 -623
rect -510 -627 -509 -623
rect -515 -629 -509 -627
rect -505 -623 -499 -621
rect -505 -627 -504 -623
rect -500 -627 -499 -623
rect -505 -629 -499 -627
rect 858 -590 864 -588
rect 868 -590 885 -582
rect 889 -584 906 -582
rect 889 -588 892 -584
rect 896 -588 906 -584
rect 889 -590 906 -588
rect 924 -584 930 -582
rect 924 -588 925 -584
rect 929 -588 930 -584
rect 924 -590 930 -588
rect 934 -584 940 -582
rect 934 -588 935 -584
rect 939 -588 940 -584
rect 1617 -584 1623 -582
rect 934 -590 940 -588
rect 1017 -587 1023 -585
rect 1017 -591 1018 -587
rect 1022 -591 1023 -587
rect 1017 -593 1023 -591
rect 1027 -587 1044 -585
rect 1027 -591 1028 -587
rect 1032 -591 1044 -587
rect 1027 -593 1044 -591
rect 1048 -587 1065 -585
rect 1048 -591 1051 -587
rect 1055 -591 1065 -587
rect 1048 -593 1065 -591
rect 1085 -587 1091 -585
rect 1085 -591 1086 -587
rect 1090 -591 1091 -587
rect 1085 -593 1091 -591
rect 1095 -587 1101 -585
rect 1095 -591 1096 -587
rect 1100 -591 1101 -587
rect 1617 -588 1618 -584
rect 1622 -588 1623 -584
rect 1095 -593 1101 -591
rect 1617 -590 1623 -588
rect 1627 -590 1644 -582
rect 1648 -584 1665 -582
rect 1648 -588 1651 -584
rect 1655 -588 1665 -584
rect 1648 -590 1665 -588
rect 1683 -584 1689 -582
rect 1683 -588 1684 -584
rect 1688 -588 1689 -584
rect 1683 -590 1689 -588
rect 1693 -584 1699 -582
rect 1693 -588 1694 -584
rect 1698 -588 1699 -584
rect 2353 -584 2359 -582
rect 1693 -590 1699 -588
rect 1776 -587 1782 -585
rect 1776 -591 1777 -587
rect 1781 -591 1782 -587
rect 1776 -593 1782 -591
rect 1786 -587 1803 -585
rect 1786 -591 1787 -587
rect 1791 -591 1803 -587
rect 1786 -593 1803 -591
rect 1807 -587 1824 -585
rect 1807 -591 1810 -587
rect 1814 -591 1824 -587
rect 1807 -593 1824 -591
rect 1844 -587 1850 -585
rect 1844 -591 1845 -587
rect 1849 -591 1850 -587
rect 1844 -593 1850 -591
rect 1854 -587 1860 -585
rect 1854 -591 1855 -587
rect 1859 -591 1860 -587
rect 2353 -588 2354 -584
rect 2358 -588 2359 -584
rect 1854 -593 1860 -591
rect 2353 -590 2359 -588
rect 2363 -590 2380 -582
rect 2384 -584 2401 -582
rect 2384 -588 2387 -584
rect 2391 -588 2401 -584
rect 2384 -590 2401 -588
rect 2419 -584 2425 -582
rect 2419 -588 2420 -584
rect 2424 -588 2425 -584
rect 2419 -590 2425 -588
rect 2429 -584 2435 -582
rect 2429 -588 2430 -584
rect 2434 -588 2435 -584
rect 2429 -590 2435 -588
rect 2512 -587 2518 -585
rect 2512 -591 2513 -587
rect 2517 -591 2518 -587
rect 2512 -593 2518 -591
rect 2522 -587 2539 -585
rect 2522 -591 2523 -587
rect 2527 -591 2539 -587
rect 2522 -593 2539 -591
rect 2543 -587 2560 -585
rect 2543 -591 2546 -587
rect 2550 -591 2560 -587
rect 2543 -593 2560 -591
rect 2580 -587 2586 -585
rect 2580 -591 2581 -587
rect 2585 -591 2586 -587
rect 2580 -593 2586 -591
rect 2590 -587 2596 -585
rect 2590 -591 2591 -587
rect 2595 -591 2596 -587
rect 2590 -593 2596 -591
rect -196 -632 -190 -630
rect -196 -636 -195 -632
rect -191 -636 -190 -632
rect -196 -638 -190 -636
rect -186 -638 -169 -630
rect -165 -632 -148 -630
rect -165 -636 -162 -632
rect -158 -636 -148 -632
rect -165 -638 -148 -636
rect -130 -632 -124 -630
rect -130 -636 -129 -632
rect -125 -636 -124 -632
rect -130 -638 -124 -636
rect -120 -632 -114 -630
rect -120 -636 -119 -632
rect -115 -636 -114 -632
rect -120 -638 -114 -636
rect 547 -635 553 -633
rect 547 -639 548 -635
rect 552 -639 553 -635
rect 547 -641 553 -639
rect 557 -641 574 -633
rect 578 -635 595 -633
rect 578 -639 581 -635
rect 585 -639 595 -635
rect 578 -641 595 -639
rect 613 -635 619 -633
rect 613 -639 614 -635
rect 618 -639 619 -635
rect 613 -641 619 -639
rect 623 -635 629 -633
rect 623 -639 624 -635
rect 628 -639 629 -635
rect 623 -641 629 -639
rect 1306 -635 1312 -633
rect 1306 -639 1307 -635
rect 1311 -639 1312 -635
rect 1306 -641 1312 -639
rect 1316 -641 1333 -633
rect 1337 -635 1354 -633
rect 1337 -639 1340 -635
rect 1344 -639 1354 -635
rect 1337 -641 1354 -639
rect 1372 -635 1378 -633
rect 1372 -639 1373 -635
rect 1377 -639 1378 -635
rect 1372 -641 1378 -639
rect 1382 -635 1388 -633
rect 1382 -639 1383 -635
rect 1387 -639 1388 -635
rect 1382 -641 1388 -639
rect 2042 -635 2048 -633
rect 2042 -639 2043 -635
rect 2047 -639 2048 -635
rect 2042 -641 2048 -639
rect 2052 -641 2069 -633
rect 2073 -635 2090 -633
rect 2073 -639 2076 -635
rect 2080 -639 2090 -635
rect 2073 -641 2090 -639
rect 2108 -635 2114 -633
rect 2108 -639 2109 -635
rect 2113 -639 2114 -635
rect 2108 -641 2114 -639
rect 2118 -635 2124 -633
rect 2118 -639 2119 -635
rect 2123 -639 2124 -635
rect 2118 -641 2124 -639
rect -581 -715 -575 -713
rect -581 -719 -580 -715
rect -576 -719 -575 -715
rect -581 -721 -575 -719
rect -571 -721 -554 -713
rect -550 -715 -533 -713
rect -550 -719 -547 -715
rect -543 -719 -533 -715
rect -550 -721 -533 -719
rect -515 -715 -509 -713
rect -515 -719 -514 -715
rect -510 -719 -509 -715
rect -515 -721 -509 -719
rect -505 -715 -499 -713
rect -505 -719 -504 -715
rect -500 -719 -499 -715
rect -505 -721 -499 -719
rect -581 -807 -575 -805
rect -581 -811 -580 -807
rect -576 -811 -575 -807
rect -581 -813 -575 -811
rect -571 -813 -554 -805
rect -550 -807 -533 -805
rect -550 -811 -547 -807
rect -543 -811 -533 -807
rect -550 -813 -533 -811
rect -515 -807 -509 -805
rect -515 -811 -514 -807
rect -510 -811 -509 -807
rect -515 -813 -509 -811
rect -505 -807 -499 -805
rect -505 -811 -504 -807
rect -500 -811 -499 -807
rect -505 -813 -499 -811
rect -124 -856 -118 -854
rect -124 -860 -123 -856
rect -119 -860 -118 -856
rect -124 -862 -118 -860
rect -114 -862 -97 -854
rect -93 -856 -76 -854
rect -93 -860 -90 -856
rect -86 -860 -76 -856
rect 474 -856 480 -854
rect -93 -862 -76 -860
rect 474 -860 475 -856
rect 479 -860 480 -856
rect 474 -862 480 -860
rect 484 -862 501 -854
rect 505 -856 522 -854
rect 505 -860 508 -856
rect 512 -860 522 -856
rect 1353 -856 1359 -854
rect 505 -862 522 -860
rect -197 -904 -191 -902
rect -197 -908 -196 -904
rect -192 -908 -191 -904
rect -197 -910 -191 -908
rect -187 -910 -170 -902
rect -166 -904 -149 -902
rect -166 -908 -163 -904
rect -159 -908 -149 -904
rect -166 -910 -149 -908
rect 1353 -860 1354 -856
rect 1358 -860 1359 -856
rect 1353 -862 1359 -860
rect 1363 -862 1380 -854
rect 1384 -856 1401 -854
rect 1384 -860 1387 -856
rect 1391 -860 1401 -856
rect 2121 -856 2127 -854
rect 1384 -862 1401 -860
rect 401 -904 407 -902
rect 401 -908 402 -904
rect 406 -908 407 -904
rect 401 -910 407 -908
rect 411 -910 428 -902
rect 432 -904 449 -902
rect 432 -908 435 -904
rect 439 -908 449 -904
rect 432 -910 449 -908
rect -23 -924 -17 -922
rect -580 -957 -574 -955
rect -580 -961 -579 -957
rect -575 -961 -574 -957
rect -580 -963 -574 -961
rect -570 -963 -553 -955
rect -549 -957 -532 -955
rect -549 -961 -546 -957
rect -542 -961 -532 -957
rect -549 -963 -532 -961
rect -514 -957 -508 -955
rect -514 -961 -513 -957
rect -509 -961 -508 -957
rect -514 -963 -508 -961
rect -504 -957 -498 -955
rect -504 -961 -503 -957
rect -499 -961 -498 -957
rect -504 -963 -498 -961
rect -23 -928 -22 -924
rect -18 -928 -17 -924
rect -23 -930 -17 -928
rect -13 -930 4 -922
rect 8 -924 25 -922
rect 8 -928 11 -924
rect 15 -928 25 -924
rect 2121 -860 2122 -856
rect 2126 -860 2127 -856
rect 2121 -862 2127 -860
rect 2131 -862 2148 -854
rect 2152 -856 2169 -854
rect 2152 -860 2155 -856
rect 2159 -860 2169 -856
rect 2152 -862 2169 -860
rect 1280 -904 1286 -902
rect 1280 -908 1281 -904
rect 1285 -908 1286 -904
rect 1280 -910 1286 -908
rect 1290 -910 1307 -902
rect 1311 -904 1328 -902
rect 1311 -908 1314 -904
rect 1318 -908 1328 -904
rect 1311 -910 1328 -908
rect 575 -924 581 -922
rect 8 -930 25 -928
rect 575 -928 576 -924
rect 580 -928 581 -924
rect 575 -930 581 -928
rect 585 -930 602 -922
rect 606 -924 623 -922
rect 606 -928 609 -924
rect 613 -928 623 -924
rect 2048 -904 2054 -902
rect 2048 -908 2049 -904
rect 2053 -908 2054 -904
rect 2048 -910 2054 -908
rect 2058 -910 2075 -902
rect 2079 -904 2096 -902
rect 2079 -908 2082 -904
rect 2086 -908 2096 -904
rect 2079 -910 2096 -908
rect 1454 -924 1460 -922
rect 606 -930 623 -928
rect 1454 -928 1455 -924
rect 1459 -928 1460 -924
rect 1454 -930 1460 -928
rect 1464 -930 1481 -922
rect 1485 -924 1502 -922
rect 1485 -928 1488 -924
rect 1492 -928 1502 -924
rect 2222 -924 2228 -922
rect 1485 -930 1502 -928
rect 2222 -928 2223 -924
rect 2227 -928 2228 -924
rect 2222 -930 2228 -928
rect 2232 -930 2249 -922
rect 2253 -924 2270 -922
rect 2253 -928 2256 -924
rect 2260 -928 2270 -924
rect 2253 -930 2270 -928
rect -109 -965 -103 -963
rect -109 -969 -108 -965
rect -104 -969 -103 -965
rect -109 -971 -103 -969
rect -99 -971 -82 -963
rect -78 -965 -61 -963
rect -78 -969 -75 -965
rect -71 -969 -61 -965
rect -78 -971 -61 -969
rect 489 -965 495 -963
rect 489 -969 490 -965
rect 494 -969 495 -965
rect 489 -971 495 -969
rect 499 -971 516 -963
rect 520 -965 537 -963
rect 520 -969 523 -965
rect 527 -969 537 -965
rect 520 -971 537 -969
rect 1368 -965 1374 -963
rect 1368 -969 1369 -965
rect 1373 -969 1374 -965
rect 1368 -971 1374 -969
rect 1378 -971 1395 -963
rect 1399 -965 1416 -963
rect 1399 -969 1402 -965
rect 1406 -969 1416 -965
rect 1399 -971 1416 -969
rect 2136 -965 2142 -963
rect 2136 -969 2137 -965
rect 2141 -969 2142 -965
rect 2136 -971 2142 -969
rect 2146 -971 2163 -963
rect 2167 -965 2184 -963
rect 2167 -969 2170 -965
rect 2174 -969 2184 -965
rect 2167 -971 2184 -969
rect -583 -1049 -577 -1047
rect -583 -1053 -582 -1049
rect -578 -1053 -577 -1049
rect -583 -1055 -577 -1053
rect -573 -1055 -556 -1047
rect -552 -1049 -535 -1047
rect -552 -1053 -549 -1049
rect -545 -1053 -535 -1049
rect -552 -1055 -535 -1053
rect -517 -1049 -511 -1047
rect -517 -1053 -516 -1049
rect -512 -1053 -511 -1049
rect -517 -1055 -511 -1053
rect -507 -1049 -501 -1047
rect -507 -1053 -506 -1049
rect -502 -1053 -501 -1049
rect -507 -1055 -501 -1053
rect -583 -1141 -577 -1139
rect -583 -1145 -582 -1141
rect -578 -1145 -577 -1141
rect -583 -1147 -577 -1145
rect -573 -1147 -556 -1139
rect -552 -1141 -535 -1139
rect -552 -1145 -549 -1141
rect -545 -1145 -535 -1141
rect -552 -1147 -535 -1145
rect -517 -1141 -511 -1139
rect -517 -1145 -516 -1141
rect -512 -1145 -511 -1141
rect -517 -1147 -511 -1145
rect -507 -1141 -501 -1139
rect -507 -1145 -506 -1141
rect -502 -1145 -501 -1141
rect -507 -1147 -501 -1145
rect 157 -1159 163 -1157
rect 157 -1163 158 -1159
rect 162 -1163 163 -1159
rect 157 -1165 163 -1163
rect 167 -1165 184 -1157
rect 188 -1159 205 -1157
rect 188 -1163 191 -1159
rect 195 -1163 205 -1159
rect 900 -1162 906 -1160
rect 188 -1165 205 -1163
rect 900 -1166 901 -1162
rect 905 -1166 906 -1162
rect 900 -1168 906 -1166
rect 910 -1168 927 -1160
rect 931 -1162 948 -1160
rect 931 -1166 934 -1162
rect 938 -1166 948 -1162
rect 1659 -1162 1665 -1160
rect 931 -1168 948 -1166
rect -153 -1207 -147 -1205
rect -153 -1211 -152 -1207
rect -148 -1211 -147 -1207
rect -153 -1213 -147 -1211
rect -143 -1213 -126 -1205
rect -122 -1207 -105 -1205
rect -122 -1211 -119 -1207
rect -115 -1211 -105 -1207
rect -122 -1213 -105 -1211
rect 84 -1207 90 -1205
rect 84 -1211 85 -1207
rect 89 -1211 90 -1207
rect 84 -1213 90 -1211
rect 94 -1213 111 -1205
rect 115 -1207 132 -1205
rect 115 -1211 118 -1207
rect 122 -1211 132 -1207
rect 115 -1213 132 -1211
rect -583 -1233 -577 -1231
rect -583 -1237 -582 -1233
rect -578 -1237 -577 -1233
rect -583 -1239 -577 -1237
rect -573 -1239 -556 -1231
rect -552 -1233 -535 -1231
rect -552 -1237 -549 -1233
rect -545 -1237 -535 -1233
rect -552 -1239 -535 -1237
rect -517 -1233 -511 -1231
rect -517 -1237 -516 -1233
rect -512 -1237 -511 -1233
rect -517 -1239 -511 -1237
rect -507 -1233 -501 -1231
rect -507 -1237 -506 -1233
rect -502 -1237 -501 -1233
rect -507 -1239 -501 -1237
rect 1659 -1166 1660 -1162
rect 1664 -1166 1665 -1162
rect 1659 -1168 1665 -1166
rect 1669 -1168 1686 -1160
rect 1690 -1162 1707 -1160
rect 1690 -1166 1693 -1162
rect 1697 -1166 1707 -1162
rect 2395 -1162 2401 -1160
rect 1690 -1168 1707 -1166
rect 590 -1210 596 -1208
rect 590 -1214 591 -1210
rect 595 -1214 596 -1210
rect 590 -1216 596 -1214
rect 600 -1216 617 -1208
rect 621 -1210 638 -1208
rect 621 -1214 624 -1210
rect 628 -1214 638 -1210
rect 621 -1216 638 -1214
rect 827 -1210 833 -1208
rect 827 -1214 828 -1210
rect 832 -1214 833 -1210
rect 827 -1216 833 -1214
rect 837 -1216 854 -1208
rect 858 -1210 875 -1208
rect 858 -1214 861 -1210
rect 865 -1214 875 -1210
rect 858 -1216 875 -1214
rect 258 -1227 264 -1225
rect -226 -1255 -220 -1253
rect -226 -1259 -225 -1255
rect -221 -1259 -220 -1255
rect -226 -1261 -220 -1259
rect -216 -1261 -199 -1253
rect -195 -1255 -178 -1253
rect -195 -1259 -192 -1255
rect -188 -1259 -178 -1255
rect -195 -1261 -178 -1259
rect 258 -1231 259 -1227
rect 263 -1231 264 -1227
rect 258 -1233 264 -1231
rect 268 -1233 285 -1225
rect 289 -1227 306 -1225
rect 289 -1231 292 -1227
rect 296 -1231 306 -1227
rect 289 -1233 306 -1231
rect 2395 -1166 2396 -1162
rect 2400 -1166 2401 -1162
rect 2395 -1168 2401 -1166
rect 2405 -1168 2422 -1160
rect 2426 -1162 2443 -1160
rect 2426 -1166 2429 -1162
rect 2433 -1166 2443 -1162
rect 2426 -1168 2443 -1166
rect 1349 -1210 1355 -1208
rect 1349 -1214 1350 -1210
rect 1354 -1214 1355 -1210
rect 1349 -1216 1355 -1214
rect 1359 -1216 1376 -1208
rect 1380 -1210 1397 -1208
rect 1380 -1214 1383 -1210
rect 1387 -1214 1397 -1210
rect 1380 -1216 1397 -1214
rect 1586 -1210 1592 -1208
rect 1586 -1214 1587 -1210
rect 1591 -1214 1592 -1210
rect 1586 -1216 1592 -1214
rect 1596 -1216 1613 -1208
rect 1617 -1210 1634 -1208
rect 1617 -1214 1620 -1210
rect 1624 -1214 1634 -1210
rect 1617 -1216 1634 -1214
rect 1001 -1230 1007 -1228
rect 517 -1258 523 -1256
rect 517 -1262 518 -1258
rect 522 -1262 523 -1258
rect 517 -1264 523 -1262
rect 527 -1264 544 -1256
rect 548 -1258 565 -1256
rect 548 -1262 551 -1258
rect 555 -1262 565 -1258
rect 548 -1264 565 -1262
rect 172 -1268 178 -1266
rect 172 -1272 173 -1268
rect 177 -1272 178 -1268
rect -52 -1275 -46 -1273
rect -52 -1279 -51 -1275
rect -47 -1279 -46 -1275
rect -52 -1281 -46 -1279
rect -42 -1281 -25 -1273
rect -21 -1275 -4 -1273
rect 172 -1274 178 -1272
rect 182 -1274 199 -1266
rect 203 -1268 220 -1266
rect 203 -1272 206 -1268
rect 210 -1272 220 -1268
rect 203 -1274 220 -1272
rect -21 -1279 -18 -1275
rect -14 -1279 -4 -1275
rect -21 -1281 -4 -1279
rect 1001 -1234 1002 -1230
rect 1006 -1234 1007 -1230
rect 1001 -1236 1007 -1234
rect 1011 -1236 1028 -1228
rect 1032 -1230 1049 -1228
rect 1032 -1234 1035 -1230
rect 1039 -1234 1049 -1230
rect 1032 -1236 1049 -1234
rect 2085 -1210 2091 -1208
rect 2085 -1214 2086 -1210
rect 2090 -1214 2091 -1210
rect 2085 -1216 2091 -1214
rect 2095 -1216 2112 -1208
rect 2116 -1210 2133 -1208
rect 2116 -1214 2119 -1210
rect 2123 -1214 2133 -1210
rect 2116 -1216 2133 -1214
rect 2322 -1210 2328 -1208
rect 2322 -1214 2323 -1210
rect 2327 -1214 2328 -1210
rect 2322 -1216 2328 -1214
rect 2332 -1216 2349 -1208
rect 2353 -1210 2370 -1208
rect 2353 -1214 2356 -1210
rect 2360 -1214 2370 -1210
rect 2353 -1216 2370 -1214
rect 1760 -1230 1766 -1228
rect 1276 -1258 1282 -1256
rect 1276 -1262 1277 -1258
rect 1281 -1262 1282 -1258
rect 1276 -1264 1282 -1262
rect 1286 -1264 1303 -1256
rect 1307 -1258 1324 -1256
rect 1307 -1262 1310 -1258
rect 1314 -1262 1324 -1258
rect 1307 -1264 1324 -1262
rect 915 -1271 921 -1269
rect 915 -1275 916 -1271
rect 920 -1275 921 -1271
rect 691 -1278 697 -1276
rect -138 -1316 -132 -1314
rect -138 -1320 -137 -1316
rect -133 -1320 -132 -1316
rect -138 -1322 -132 -1320
rect -128 -1322 -111 -1314
rect -107 -1316 -90 -1314
rect -107 -1320 -104 -1316
rect -100 -1320 -90 -1316
rect 691 -1282 692 -1278
rect 696 -1282 697 -1278
rect 691 -1284 697 -1282
rect 701 -1284 718 -1276
rect 722 -1278 739 -1276
rect 915 -1277 921 -1275
rect 925 -1277 942 -1269
rect 946 -1271 963 -1269
rect 946 -1275 949 -1271
rect 953 -1275 963 -1271
rect 946 -1277 963 -1275
rect 722 -1282 725 -1278
rect 729 -1282 739 -1278
rect 722 -1284 739 -1282
rect 1760 -1234 1761 -1230
rect 1765 -1234 1766 -1230
rect 1760 -1236 1766 -1234
rect 1770 -1236 1787 -1228
rect 1791 -1230 1808 -1228
rect 1791 -1234 1794 -1230
rect 1798 -1234 1808 -1230
rect 1791 -1236 1808 -1234
rect 2496 -1230 2502 -1228
rect 2012 -1258 2018 -1256
rect 2012 -1262 2013 -1258
rect 2017 -1262 2018 -1258
rect 2012 -1264 2018 -1262
rect 2022 -1264 2039 -1256
rect 2043 -1258 2060 -1256
rect 2043 -1262 2046 -1258
rect 2050 -1262 2060 -1258
rect 2043 -1264 2060 -1262
rect 1674 -1271 1680 -1269
rect 1674 -1275 1675 -1271
rect 1679 -1275 1680 -1271
rect 1450 -1278 1456 -1276
rect 1450 -1282 1451 -1278
rect 1455 -1282 1456 -1278
rect 1450 -1284 1456 -1282
rect 1460 -1284 1477 -1276
rect 1481 -1278 1498 -1276
rect 1674 -1277 1680 -1275
rect 1684 -1277 1701 -1269
rect 1705 -1271 1722 -1269
rect 1705 -1275 1708 -1271
rect 1712 -1275 1722 -1271
rect 1705 -1277 1722 -1275
rect 1481 -1282 1484 -1278
rect 1488 -1282 1498 -1278
rect 1481 -1284 1498 -1282
rect 2496 -1234 2497 -1230
rect 2501 -1234 2502 -1230
rect 2496 -1236 2502 -1234
rect 2506 -1236 2523 -1228
rect 2527 -1230 2544 -1228
rect 2527 -1234 2530 -1230
rect 2534 -1234 2544 -1230
rect 2527 -1236 2544 -1234
rect 2410 -1271 2416 -1269
rect 2410 -1275 2411 -1271
rect 2415 -1275 2416 -1271
rect 2186 -1278 2192 -1276
rect 2186 -1282 2187 -1278
rect 2191 -1282 2192 -1278
rect 2186 -1284 2192 -1282
rect 2196 -1284 2213 -1276
rect 2217 -1278 2234 -1276
rect 2410 -1277 2416 -1275
rect 2420 -1277 2437 -1269
rect 2441 -1271 2458 -1269
rect 2441 -1275 2444 -1271
rect 2448 -1275 2458 -1271
rect 2441 -1277 2458 -1275
rect 2217 -1282 2220 -1278
rect 2224 -1282 2234 -1278
rect 2217 -1284 2234 -1282
rect -107 -1322 -90 -1320
rect 605 -1319 611 -1317
rect -578 -1324 -572 -1322
rect -578 -1328 -577 -1324
rect -573 -1328 -572 -1324
rect -578 -1330 -572 -1328
rect -568 -1330 -551 -1322
rect -547 -1324 -530 -1322
rect -547 -1328 -544 -1324
rect -540 -1328 -530 -1324
rect -547 -1330 -530 -1328
rect -512 -1324 -506 -1322
rect -512 -1328 -511 -1324
rect -507 -1328 -506 -1324
rect -512 -1330 -506 -1328
rect -502 -1324 -496 -1322
rect -502 -1328 -501 -1324
rect -497 -1328 -496 -1324
rect -502 -1330 -496 -1328
rect 605 -1323 606 -1319
rect 610 -1323 611 -1319
rect 605 -1325 611 -1323
rect 615 -1325 632 -1317
rect 636 -1319 653 -1317
rect 636 -1323 639 -1319
rect 643 -1323 653 -1319
rect 636 -1325 653 -1323
rect 1364 -1319 1370 -1317
rect 1364 -1323 1365 -1319
rect 1369 -1323 1370 -1319
rect 1364 -1325 1370 -1323
rect 1374 -1325 1391 -1317
rect 1395 -1319 1412 -1317
rect 1395 -1323 1398 -1319
rect 1402 -1323 1412 -1319
rect 1395 -1325 1412 -1323
rect 2100 -1319 2106 -1317
rect 2100 -1323 2101 -1319
rect 2105 -1323 2106 -1319
rect 2100 -1325 2106 -1323
rect 2110 -1325 2127 -1317
rect 2131 -1319 2148 -1317
rect 2131 -1323 2134 -1319
rect 2138 -1323 2148 -1319
rect 2131 -1325 2148 -1323
rect 144 -1374 150 -1372
rect 144 -1378 145 -1374
rect 149 -1378 150 -1374
rect 144 -1380 150 -1378
rect 154 -1380 171 -1372
rect 175 -1374 192 -1372
rect 175 -1378 178 -1374
rect 182 -1378 192 -1374
rect 175 -1380 192 -1378
rect 210 -1374 216 -1372
rect 210 -1378 211 -1374
rect 215 -1378 216 -1374
rect 210 -1380 216 -1378
rect 220 -1374 226 -1372
rect 220 -1378 221 -1374
rect 225 -1378 226 -1374
rect 220 -1380 226 -1378
rect 303 -1377 309 -1375
rect 303 -1381 304 -1377
rect 308 -1381 309 -1377
rect 303 -1383 309 -1381
rect 313 -1377 330 -1375
rect 313 -1381 314 -1377
rect 318 -1381 330 -1377
rect 313 -1383 330 -1381
rect 334 -1377 351 -1375
rect 334 -1381 337 -1377
rect 341 -1381 351 -1377
rect 334 -1383 351 -1381
rect 371 -1377 377 -1375
rect 371 -1381 372 -1377
rect 376 -1381 377 -1377
rect 371 -1383 377 -1381
rect 381 -1377 387 -1375
rect 381 -1381 382 -1377
rect 386 -1381 387 -1377
rect 887 -1377 893 -1375
rect 887 -1381 888 -1377
rect 892 -1381 893 -1377
rect 381 -1383 387 -1381
rect -581 -1416 -575 -1414
rect -581 -1420 -580 -1416
rect -576 -1420 -575 -1416
rect -581 -1422 -575 -1420
rect -571 -1422 -554 -1414
rect -550 -1416 -533 -1414
rect -550 -1420 -547 -1416
rect -543 -1420 -533 -1416
rect -550 -1422 -533 -1420
rect -515 -1416 -509 -1414
rect -515 -1420 -514 -1416
rect -510 -1420 -509 -1416
rect -515 -1422 -509 -1420
rect -505 -1416 -499 -1414
rect -505 -1420 -504 -1416
rect -500 -1420 -499 -1416
rect -505 -1422 -499 -1420
rect 887 -1383 893 -1381
rect 897 -1383 914 -1375
rect 918 -1377 935 -1375
rect 918 -1381 921 -1377
rect 925 -1381 935 -1377
rect 918 -1383 935 -1381
rect 953 -1377 959 -1375
rect 953 -1381 954 -1377
rect 958 -1381 959 -1377
rect 953 -1383 959 -1381
rect 963 -1377 969 -1375
rect 963 -1381 964 -1377
rect 968 -1381 969 -1377
rect 1646 -1377 1652 -1375
rect 963 -1383 969 -1381
rect 1046 -1380 1052 -1378
rect 1046 -1384 1047 -1380
rect 1051 -1384 1052 -1380
rect 1046 -1386 1052 -1384
rect 1056 -1380 1073 -1378
rect 1056 -1384 1057 -1380
rect 1061 -1384 1073 -1380
rect 1056 -1386 1073 -1384
rect 1077 -1380 1094 -1378
rect 1077 -1384 1080 -1380
rect 1084 -1384 1094 -1380
rect 1077 -1386 1094 -1384
rect 1114 -1380 1120 -1378
rect 1114 -1384 1115 -1380
rect 1119 -1384 1120 -1380
rect 1114 -1386 1120 -1384
rect 1124 -1380 1130 -1378
rect 1124 -1384 1125 -1380
rect 1129 -1384 1130 -1380
rect 1646 -1381 1647 -1377
rect 1651 -1381 1652 -1377
rect 1124 -1386 1130 -1384
rect 1646 -1383 1652 -1381
rect 1656 -1383 1673 -1375
rect 1677 -1377 1694 -1375
rect 1677 -1381 1680 -1377
rect 1684 -1381 1694 -1377
rect 1677 -1383 1694 -1381
rect 1712 -1377 1718 -1375
rect 1712 -1381 1713 -1377
rect 1717 -1381 1718 -1377
rect 1712 -1383 1718 -1381
rect 1722 -1377 1728 -1375
rect 1722 -1381 1723 -1377
rect 1727 -1381 1728 -1377
rect 2382 -1377 2388 -1375
rect 1722 -1383 1728 -1381
rect 1805 -1380 1811 -1378
rect 1805 -1384 1806 -1380
rect 1810 -1384 1811 -1380
rect 1805 -1386 1811 -1384
rect 1815 -1380 1832 -1378
rect 1815 -1384 1816 -1380
rect 1820 -1384 1832 -1380
rect 1815 -1386 1832 -1384
rect 1836 -1380 1853 -1378
rect 1836 -1384 1839 -1380
rect 1843 -1384 1853 -1380
rect 1836 -1386 1853 -1384
rect 1873 -1380 1879 -1378
rect 1873 -1384 1874 -1380
rect 1878 -1384 1879 -1380
rect 1873 -1386 1879 -1384
rect 1883 -1380 1889 -1378
rect 1883 -1384 1884 -1380
rect 1888 -1384 1889 -1380
rect 2382 -1381 2383 -1377
rect 2387 -1381 2388 -1377
rect 1883 -1386 1889 -1384
rect 2382 -1383 2388 -1381
rect 2392 -1383 2409 -1375
rect 2413 -1377 2430 -1375
rect 2413 -1381 2416 -1377
rect 2420 -1381 2430 -1377
rect 2413 -1383 2430 -1381
rect 2448 -1377 2454 -1375
rect 2448 -1381 2449 -1377
rect 2453 -1381 2454 -1377
rect 2448 -1383 2454 -1381
rect 2458 -1377 2464 -1375
rect 2458 -1381 2459 -1377
rect 2463 -1381 2464 -1377
rect 2458 -1383 2464 -1381
rect 2541 -1380 2547 -1378
rect 2541 -1384 2542 -1380
rect 2546 -1384 2547 -1380
rect 2541 -1386 2547 -1384
rect 2551 -1380 2568 -1378
rect 2551 -1384 2552 -1380
rect 2556 -1384 2568 -1380
rect 2551 -1386 2568 -1384
rect 2572 -1380 2589 -1378
rect 2572 -1384 2575 -1380
rect 2579 -1384 2589 -1380
rect 2572 -1386 2589 -1384
rect 2609 -1380 2615 -1378
rect 2609 -1384 2610 -1380
rect 2614 -1384 2615 -1380
rect 2609 -1386 2615 -1384
rect 2619 -1380 2625 -1378
rect 2619 -1384 2620 -1380
rect 2624 -1384 2625 -1380
rect 2619 -1386 2625 -1384
rect -167 -1425 -161 -1423
rect -167 -1429 -166 -1425
rect -162 -1429 -161 -1425
rect -167 -1431 -161 -1429
rect -157 -1431 -140 -1423
rect -136 -1425 -119 -1423
rect -136 -1429 -133 -1425
rect -129 -1429 -119 -1425
rect -136 -1431 -119 -1429
rect -101 -1425 -95 -1423
rect -101 -1429 -100 -1425
rect -96 -1429 -95 -1425
rect -101 -1431 -95 -1429
rect -91 -1425 -85 -1423
rect -91 -1429 -90 -1425
rect -86 -1429 -85 -1425
rect -91 -1431 -85 -1429
rect 576 -1428 582 -1426
rect 576 -1432 577 -1428
rect 581 -1432 582 -1428
rect 576 -1434 582 -1432
rect 586 -1434 603 -1426
rect 607 -1428 624 -1426
rect 607 -1432 610 -1428
rect 614 -1432 624 -1428
rect 607 -1434 624 -1432
rect 642 -1428 648 -1426
rect 642 -1432 643 -1428
rect 647 -1432 648 -1428
rect 642 -1434 648 -1432
rect 652 -1428 658 -1426
rect 652 -1432 653 -1428
rect 657 -1432 658 -1428
rect 652 -1434 658 -1432
rect 1335 -1428 1341 -1426
rect 1335 -1432 1336 -1428
rect 1340 -1432 1341 -1428
rect 1335 -1434 1341 -1432
rect 1345 -1434 1362 -1426
rect 1366 -1428 1383 -1426
rect 1366 -1432 1369 -1428
rect 1373 -1432 1383 -1428
rect 1366 -1434 1383 -1432
rect 1401 -1428 1407 -1426
rect 1401 -1432 1402 -1428
rect 1406 -1432 1407 -1428
rect 1401 -1434 1407 -1432
rect 1411 -1428 1417 -1426
rect 1411 -1432 1412 -1428
rect 1416 -1432 1417 -1428
rect 1411 -1434 1417 -1432
rect 2071 -1428 2077 -1426
rect 2071 -1432 2072 -1428
rect 2076 -1432 2077 -1428
rect 2071 -1434 2077 -1432
rect 2081 -1434 2098 -1426
rect 2102 -1428 2119 -1426
rect 2102 -1432 2105 -1428
rect 2109 -1432 2119 -1428
rect 2102 -1434 2119 -1432
rect 2137 -1428 2143 -1426
rect 2137 -1432 2138 -1428
rect 2142 -1432 2143 -1428
rect 2137 -1434 2143 -1432
rect 2147 -1428 2153 -1426
rect 2147 -1432 2148 -1428
rect 2152 -1432 2153 -1428
rect 2147 -1434 2153 -1432
rect -581 -1508 -575 -1506
rect -581 -1512 -580 -1508
rect -576 -1512 -575 -1508
rect -581 -1514 -575 -1512
rect -571 -1514 -554 -1506
rect -550 -1508 -533 -1506
rect -550 -1512 -547 -1508
rect -543 -1512 -533 -1508
rect -550 -1514 -533 -1512
rect -515 -1508 -509 -1506
rect -515 -1512 -514 -1508
rect -510 -1512 -509 -1508
rect -515 -1514 -509 -1512
rect -505 -1508 -499 -1506
rect -505 -1512 -504 -1508
rect -500 -1512 -499 -1508
rect -505 -1514 -499 -1512
rect -581 -1600 -575 -1598
rect -581 -1604 -580 -1600
rect -576 -1604 -575 -1600
rect -581 -1606 -575 -1604
rect -571 -1606 -554 -1598
rect -550 -1600 -533 -1598
rect -550 -1604 -547 -1600
rect -543 -1604 -533 -1600
rect -550 -1606 -533 -1604
rect -515 -1600 -509 -1598
rect -515 -1604 -514 -1600
rect -510 -1604 -509 -1600
rect -515 -1606 -509 -1604
rect -505 -1600 -499 -1598
rect -505 -1604 -504 -1600
rect -500 -1604 -499 -1600
rect -505 -1606 -499 -1604
rect -580 -1720 -574 -1718
rect -580 -1724 -579 -1720
rect -575 -1724 -574 -1720
rect -580 -1726 -574 -1724
rect -570 -1726 -553 -1718
rect -549 -1720 -532 -1718
rect -549 -1724 -546 -1720
rect -542 -1724 -532 -1720
rect -549 -1726 -532 -1724
rect -514 -1720 -508 -1718
rect -514 -1724 -513 -1720
rect -509 -1724 -508 -1720
rect -514 -1726 -508 -1724
rect -504 -1720 -498 -1718
rect -504 -1724 -503 -1720
rect -499 -1724 -498 -1720
rect -504 -1726 -498 -1724
rect 13 -1776 19 -1774
rect 13 -1780 14 -1776
rect 18 -1780 19 -1776
rect 13 -1782 19 -1780
rect 23 -1782 40 -1774
rect 44 -1776 61 -1774
rect 44 -1780 47 -1776
rect 51 -1780 61 -1776
rect 502 -1776 508 -1774
rect 44 -1782 61 -1780
rect -583 -1812 -577 -1810
rect -583 -1816 -582 -1812
rect -578 -1816 -577 -1812
rect -583 -1818 -577 -1816
rect -573 -1818 -556 -1810
rect -552 -1812 -535 -1810
rect -552 -1816 -549 -1812
rect -545 -1816 -535 -1812
rect -552 -1818 -535 -1816
rect -517 -1812 -511 -1810
rect -517 -1816 -516 -1812
rect -512 -1816 -511 -1812
rect -517 -1818 -511 -1816
rect -507 -1812 -501 -1810
rect -507 -1816 -506 -1812
rect -502 -1816 -501 -1812
rect -507 -1818 -501 -1816
rect 502 -1780 503 -1776
rect 507 -1780 508 -1776
rect 502 -1782 508 -1780
rect 512 -1782 529 -1774
rect 533 -1776 550 -1774
rect 533 -1780 536 -1776
rect 540 -1780 550 -1776
rect 886 -1776 892 -1774
rect 533 -1782 550 -1780
rect -60 -1824 -54 -1822
rect -60 -1828 -59 -1824
rect -55 -1828 -54 -1824
rect -60 -1830 -54 -1828
rect -50 -1830 -33 -1822
rect -29 -1824 -12 -1822
rect -29 -1828 -26 -1824
rect -22 -1828 -12 -1824
rect -29 -1830 -12 -1828
rect -101 -1846 -96 -1841
rect 886 -1780 887 -1776
rect 891 -1780 892 -1776
rect 886 -1782 892 -1780
rect 896 -1782 913 -1774
rect 917 -1776 934 -1774
rect 917 -1780 920 -1776
rect 924 -1780 934 -1776
rect 917 -1782 934 -1780
rect 429 -1824 435 -1822
rect 429 -1828 430 -1824
rect 434 -1828 435 -1824
rect 429 -1830 435 -1828
rect 439 -1830 456 -1822
rect 460 -1824 477 -1822
rect 460 -1828 463 -1824
rect 467 -1828 477 -1824
rect 460 -1830 477 -1828
rect 240 -1842 246 -1840
rect 114 -1844 120 -1842
rect 114 -1848 115 -1844
rect 119 -1848 120 -1844
rect 114 -1850 120 -1848
rect 124 -1850 141 -1842
rect 145 -1844 162 -1842
rect 145 -1848 148 -1844
rect 152 -1848 162 -1844
rect 240 -1846 241 -1842
rect 245 -1846 246 -1842
rect 240 -1848 246 -1846
rect 250 -1842 256 -1840
rect 250 -1846 251 -1842
rect 255 -1846 256 -1842
rect 1301 -1800 1307 -1798
rect 813 -1824 819 -1822
rect 813 -1828 814 -1824
rect 818 -1828 819 -1824
rect 813 -1830 819 -1828
rect 823 -1830 840 -1822
rect 844 -1824 861 -1822
rect 844 -1828 847 -1824
rect 851 -1828 861 -1824
rect 844 -1830 861 -1828
rect 676 -1842 682 -1840
rect 603 -1844 609 -1842
rect 250 -1848 256 -1846
rect 145 -1850 162 -1848
rect 603 -1848 604 -1844
rect 608 -1848 609 -1844
rect 603 -1850 609 -1848
rect 613 -1850 630 -1842
rect 634 -1844 651 -1842
rect 634 -1848 637 -1844
rect 641 -1848 651 -1844
rect 676 -1846 677 -1842
rect 681 -1846 682 -1842
rect 676 -1848 682 -1846
rect 686 -1842 692 -1840
rect 686 -1846 687 -1842
rect 691 -1846 692 -1842
rect 1301 -1804 1302 -1800
rect 1306 -1804 1307 -1800
rect 1301 -1806 1307 -1804
rect 1311 -1806 1328 -1798
rect 1332 -1800 1349 -1798
rect 1332 -1804 1335 -1800
rect 1339 -1804 1349 -1800
rect 1332 -1806 1349 -1804
rect 1094 -1842 1100 -1840
rect 1021 -1844 1027 -1842
rect 686 -1848 692 -1846
rect 634 -1850 651 -1848
rect 1021 -1848 1022 -1844
rect 1026 -1848 1027 -1844
rect 1021 -1850 1027 -1848
rect 1031 -1850 1048 -1842
rect 1052 -1844 1069 -1842
rect 1052 -1848 1055 -1844
rect 1059 -1848 1069 -1844
rect 1094 -1846 1095 -1842
rect 1099 -1846 1100 -1842
rect 1094 -1848 1100 -1846
rect 1104 -1842 1110 -1840
rect 1104 -1846 1105 -1842
rect 1109 -1846 1110 -1842
rect 1104 -1848 1110 -1846
rect 1228 -1848 1234 -1846
rect 1052 -1850 1069 -1848
rect 1228 -1852 1229 -1848
rect 1233 -1852 1234 -1848
rect 1228 -1854 1234 -1852
rect 1238 -1854 1255 -1846
rect 1259 -1848 1276 -1846
rect 1259 -1852 1262 -1848
rect 1266 -1852 1276 -1848
rect 1259 -1854 1276 -1852
rect 1470 -1862 1476 -1860
rect 1470 -1866 1471 -1862
rect 1475 -1866 1476 -1862
rect 1402 -1868 1408 -1866
rect 28 -1885 34 -1883
rect 28 -1889 29 -1885
rect 33 -1889 34 -1885
rect 28 -1891 34 -1889
rect 38 -1891 55 -1883
rect 59 -1885 76 -1883
rect 59 -1889 62 -1885
rect 66 -1889 76 -1885
rect 59 -1891 76 -1889
rect 517 -1885 523 -1883
rect 517 -1889 518 -1885
rect 522 -1889 523 -1885
rect 517 -1891 523 -1889
rect 527 -1891 544 -1883
rect 548 -1885 565 -1883
rect 548 -1889 551 -1885
rect 555 -1889 565 -1885
rect 548 -1891 565 -1889
rect 901 -1885 907 -1883
rect 901 -1889 902 -1885
rect 906 -1889 907 -1885
rect 901 -1891 907 -1889
rect 911 -1891 928 -1883
rect 932 -1885 949 -1883
rect 932 -1889 935 -1885
rect 939 -1889 949 -1885
rect 932 -1891 949 -1889
rect -583 -1904 -577 -1902
rect -583 -1908 -582 -1904
rect -578 -1908 -577 -1904
rect -583 -1910 -577 -1908
rect -573 -1910 -556 -1902
rect -552 -1904 -535 -1902
rect -552 -1908 -549 -1904
rect -545 -1908 -535 -1904
rect -552 -1910 -535 -1908
rect -517 -1904 -511 -1902
rect -517 -1908 -516 -1904
rect -512 -1908 -511 -1904
rect -517 -1910 -511 -1908
rect -507 -1904 -501 -1902
rect -119 -1904 -103 -1896
rect -507 -1908 -506 -1904
rect -502 -1908 -501 -1904
rect 1402 -1872 1403 -1868
rect 1407 -1872 1408 -1868
rect 1402 -1874 1408 -1872
rect 1412 -1874 1429 -1866
rect 1433 -1868 1450 -1866
rect 1470 -1868 1476 -1866
rect 1480 -1862 1486 -1860
rect 1480 -1866 1481 -1862
rect 1485 -1866 1486 -1862
rect 1480 -1868 1486 -1866
rect 1433 -1872 1436 -1868
rect 1440 -1872 1450 -1868
rect 1433 -1874 1450 -1872
rect -507 -1910 -501 -1908
rect 1316 -1909 1322 -1907
rect 1316 -1913 1317 -1909
rect 1321 -1913 1322 -1909
rect 1316 -1915 1322 -1913
rect 1326 -1915 1343 -1907
rect 1347 -1909 1364 -1907
rect 1347 -1913 1350 -1909
rect 1354 -1913 1364 -1909
rect 1347 -1915 1364 -1913
rect -583 -1996 -577 -1994
rect -583 -2000 -582 -1996
rect -578 -2000 -577 -1996
rect -583 -2002 -577 -2000
rect -573 -2002 -556 -1994
rect -552 -1996 -535 -1994
rect -552 -2000 -549 -1996
rect -545 -2000 -535 -1996
rect -552 -2002 -535 -2000
rect -517 -1996 -511 -1994
rect -517 -2000 -516 -1996
rect -512 -2000 -511 -1996
rect -517 -2002 -511 -2000
rect -507 -1996 -501 -1994
rect -507 -2000 -506 -1996
rect -502 -2000 -501 -1996
rect -507 -2002 -501 -2000
rect -170 -2004 -165 -1996
rect -202 -2021 -197 -2013
rect -213 -2046 -208 -2038
rect -578 -2087 -572 -2085
rect -578 -2091 -577 -2087
rect -573 -2091 -572 -2087
rect -578 -2093 -572 -2091
rect -568 -2093 -551 -2085
rect -547 -2087 -530 -2085
rect -547 -2091 -544 -2087
rect -540 -2091 -530 -2087
rect -547 -2093 -530 -2091
rect -512 -2087 -506 -2085
rect -512 -2091 -511 -2087
rect -507 -2091 -506 -2087
rect -512 -2093 -506 -2091
rect -502 -2087 -496 -2085
rect -502 -2091 -501 -2087
rect -497 -2091 -496 -2087
rect -502 -2093 -496 -2091
rect -581 -2179 -575 -2177
rect -581 -2183 -580 -2179
rect -576 -2183 -575 -2179
rect -581 -2185 -575 -2183
rect -571 -2185 -554 -2177
rect -550 -2179 -533 -2177
rect -550 -2183 -547 -2179
rect -543 -2183 -533 -2179
rect -550 -2185 -533 -2183
rect -515 -2179 -509 -2177
rect -515 -2183 -514 -2179
rect -510 -2183 -509 -2179
rect -515 -2185 -509 -2183
rect -505 -2179 -499 -2177
rect -505 -2183 -504 -2179
rect -500 -2183 -499 -2179
rect -505 -2185 -499 -2183
rect -34 -2205 -28 -2203
rect -34 -2209 -33 -2205
rect -29 -2209 -28 -2205
rect -34 -2211 -28 -2209
rect -24 -2205 -18 -2203
rect -24 -2209 -23 -2205
rect -19 -2209 -18 -2205
rect -24 -2211 -18 -2209
rect 333 -2163 339 -2161
rect 333 -2167 334 -2163
rect 338 -2167 339 -2163
rect 333 -2169 339 -2167
rect 343 -2169 372 -2161
rect 376 -2169 396 -2161
rect 400 -2163 418 -2161
rect 400 -2167 407 -2163
rect 411 -2167 418 -2163
rect 400 -2169 418 -2167
rect 441 -2163 447 -2161
rect 441 -2167 442 -2163
rect 446 -2167 447 -2163
rect 441 -2169 447 -2167
rect 451 -2163 457 -2161
rect 451 -2167 452 -2163
rect 456 -2167 457 -2163
rect 451 -2169 457 -2167
rect 749 -2163 755 -2161
rect 749 -2167 750 -2163
rect 754 -2167 755 -2163
rect 749 -2169 755 -2167
rect 759 -2169 788 -2161
rect 792 -2169 812 -2161
rect 816 -2163 834 -2161
rect 816 -2167 823 -2163
rect 827 -2167 834 -2163
rect 816 -2169 834 -2167
rect 857 -2163 863 -2161
rect 857 -2167 858 -2163
rect 862 -2167 863 -2163
rect 857 -2169 863 -2167
rect 867 -2163 873 -2161
rect 867 -2167 868 -2163
rect 872 -2167 873 -2163
rect 867 -2169 873 -2167
rect 1199 -2163 1205 -2161
rect 1199 -2167 1200 -2163
rect 1204 -2167 1205 -2163
rect 1199 -2169 1205 -2167
rect 1209 -2169 1238 -2161
rect 1242 -2169 1262 -2161
rect 1266 -2163 1284 -2161
rect 1266 -2167 1273 -2163
rect 1277 -2167 1284 -2163
rect 1266 -2169 1284 -2167
rect 1307 -2163 1313 -2161
rect 1307 -2167 1308 -2163
rect 1312 -2167 1313 -2163
rect 1307 -2169 1313 -2167
rect 1317 -2163 1323 -2161
rect 1317 -2167 1318 -2163
rect 1322 -2167 1323 -2163
rect 1317 -2169 1323 -2167
rect 255 -2187 261 -2185
rect 255 -2191 256 -2187
rect 260 -2191 261 -2187
rect 255 -2193 261 -2191
rect 265 -2187 271 -2185
rect 265 -2191 266 -2187
rect 270 -2191 271 -2187
rect 265 -2193 271 -2191
rect 671 -2187 677 -2185
rect 671 -2191 672 -2187
rect 676 -2191 677 -2187
rect 671 -2193 677 -2191
rect 681 -2187 687 -2185
rect 681 -2191 682 -2187
rect 686 -2191 687 -2187
rect 681 -2193 687 -2191
rect 1115 -2187 1121 -2185
rect 1115 -2191 1116 -2187
rect 1120 -2191 1121 -2187
rect 1115 -2193 1121 -2191
rect 1125 -2187 1131 -2185
rect 1125 -2191 1126 -2187
rect 1130 -2191 1131 -2187
rect 1125 -2193 1131 -2191
rect 195 -2208 200 -2203
rect 1052 -2208 1057 -2203
rect 53 -2219 59 -2217
rect 53 -2223 54 -2219
rect 58 -2223 59 -2219
rect 53 -2225 59 -2223
rect 63 -2225 80 -2217
rect 84 -2219 101 -2217
rect 84 -2223 87 -2219
rect 91 -2223 101 -2219
rect 84 -2225 101 -2223
rect 119 -2219 125 -2217
rect 119 -2223 120 -2219
rect 124 -2223 125 -2219
rect 119 -2225 125 -2223
rect 129 -2219 135 -2217
rect 129 -2223 130 -2219
rect 134 -2223 135 -2219
rect 129 -2225 135 -2223
rect -581 -2271 -575 -2269
rect -581 -2275 -580 -2271
rect -576 -2275 -575 -2271
rect -581 -2277 -575 -2275
rect -571 -2277 -554 -2269
rect -550 -2271 -533 -2269
rect -550 -2275 -547 -2271
rect -543 -2275 -533 -2271
rect -550 -2277 -533 -2275
rect -515 -2271 -509 -2269
rect -515 -2275 -514 -2271
rect -510 -2275 -509 -2271
rect -515 -2277 -509 -2275
rect -505 -2271 -499 -2269
rect -505 -2275 -504 -2271
rect -500 -2275 -499 -2271
rect -505 -2277 -499 -2275
rect 255 -2279 261 -2277
rect 255 -2283 256 -2279
rect 260 -2283 261 -2279
rect 255 -2285 261 -2283
rect 265 -2279 271 -2277
rect 265 -2283 266 -2279
rect 270 -2283 271 -2279
rect 265 -2285 271 -2283
rect -36 -2298 -30 -2296
rect -36 -2302 -35 -2298
rect -31 -2302 -30 -2298
rect -36 -2304 -30 -2302
rect -26 -2298 -20 -2296
rect -26 -2302 -25 -2298
rect -21 -2302 -20 -2298
rect -26 -2304 -20 -2302
rect 36 -2329 41 -2324
rect 608 -2236 613 -2231
rect 351 -2300 357 -2298
rect 351 -2304 352 -2300
rect 356 -2304 357 -2300
rect 351 -2306 357 -2304
rect 361 -2306 390 -2298
rect 394 -2306 414 -2298
rect 418 -2300 436 -2298
rect 418 -2304 425 -2300
rect 429 -2304 436 -2300
rect 418 -2306 436 -2304
rect 459 -2300 465 -2298
rect 459 -2304 460 -2300
rect 464 -2304 465 -2300
rect 459 -2306 465 -2304
rect 469 -2300 475 -2298
rect 469 -2304 470 -2300
rect 474 -2304 475 -2300
rect 469 -2306 475 -2304
rect 664 -2307 670 -2305
rect 664 -2311 665 -2307
rect 669 -2311 670 -2307
rect 664 -2313 670 -2311
rect 674 -2307 680 -2305
rect 674 -2311 675 -2307
rect 679 -2311 680 -2307
rect 674 -2313 680 -2311
rect 54 -2335 60 -2333
rect 54 -2339 55 -2335
rect 59 -2339 60 -2335
rect 54 -2341 60 -2339
rect 64 -2341 81 -2333
rect 85 -2335 102 -2333
rect 85 -2339 88 -2335
rect 92 -2339 102 -2335
rect 85 -2341 102 -2339
rect 120 -2335 126 -2333
rect 120 -2339 121 -2335
rect 125 -2339 126 -2335
rect 120 -2341 126 -2339
rect 130 -2335 136 -2333
rect 130 -2339 131 -2335
rect 135 -2339 136 -2335
rect 130 -2341 136 -2339
rect 1114 -2279 1120 -2277
rect 1114 -2283 1115 -2279
rect 1119 -2283 1120 -2279
rect 1114 -2285 1120 -2283
rect 1124 -2279 1130 -2277
rect 1124 -2283 1125 -2279
rect 1129 -2283 1130 -2279
rect 1124 -2285 1130 -2283
rect 1217 -2300 1223 -2298
rect 1217 -2304 1218 -2300
rect 1222 -2304 1223 -2300
rect 1217 -2306 1223 -2304
rect 1227 -2306 1256 -2298
rect 1260 -2306 1280 -2298
rect 1284 -2300 1302 -2298
rect 1284 -2304 1291 -2300
rect 1295 -2304 1302 -2300
rect 1284 -2306 1302 -2304
rect 1325 -2300 1331 -2298
rect 1325 -2304 1326 -2300
rect 1330 -2304 1331 -2300
rect 1325 -2306 1331 -2304
rect 1335 -2300 1341 -2298
rect 1335 -2304 1336 -2300
rect 1340 -2304 1341 -2300
rect 1335 -2306 1341 -2304
rect 956 -2317 962 -2315
rect 956 -2321 957 -2317
rect 961 -2321 962 -2317
rect 956 -2323 962 -2321
rect 966 -2323 983 -2315
rect 987 -2317 1004 -2315
rect 987 -2321 990 -2317
rect 994 -2321 1004 -2317
rect 987 -2323 1004 -2321
rect 1022 -2317 1028 -2315
rect 1022 -2321 1023 -2317
rect 1027 -2321 1028 -2317
rect 1022 -2323 1028 -2321
rect 1032 -2317 1038 -2315
rect 1032 -2321 1033 -2317
rect 1037 -2321 1038 -2317
rect 1032 -2323 1038 -2321
rect 767 -2328 773 -2326
rect 767 -2332 768 -2328
rect 772 -2332 773 -2328
rect 767 -2334 773 -2332
rect 777 -2334 806 -2326
rect 810 -2334 830 -2326
rect 834 -2328 852 -2326
rect 834 -2332 841 -2328
rect 845 -2332 852 -2328
rect 834 -2334 852 -2332
rect 875 -2328 881 -2326
rect 875 -2332 876 -2328
rect 880 -2332 881 -2328
rect 875 -2334 881 -2332
rect 885 -2328 891 -2326
rect 885 -2332 886 -2328
rect 890 -2332 891 -2328
rect 885 -2334 891 -2332
rect 1437 -2329 1443 -2327
rect 1437 -2333 1438 -2329
rect 1442 -2333 1443 -2329
rect 1437 -2335 1443 -2333
rect 1447 -2335 1472 -2327
rect 1476 -2335 1496 -2327
rect 1500 -2335 1520 -2327
rect 1524 -2329 1541 -2327
rect 1524 -2333 1530 -2329
rect 1534 -2333 1541 -2329
rect 1524 -2335 1541 -2333
rect 1561 -2329 1567 -2327
rect 1561 -2333 1562 -2329
rect 1566 -2333 1567 -2329
rect 1561 -2335 1567 -2333
rect 1571 -2329 1577 -2327
rect 1571 -2333 1572 -2329
rect 1576 -2333 1577 -2329
rect 1571 -2335 1577 -2333
rect 547 -2356 553 -2354
rect 547 -2360 548 -2356
rect 552 -2360 553 -2356
rect -581 -2363 -575 -2361
rect -581 -2367 -580 -2363
rect -576 -2367 -575 -2363
rect -581 -2369 -575 -2367
rect -571 -2369 -554 -2361
rect -550 -2363 -533 -2361
rect -550 -2367 -547 -2363
rect -543 -2367 -533 -2363
rect -550 -2369 -533 -2367
rect -515 -2363 -509 -2361
rect -515 -2367 -514 -2363
rect -510 -2367 -509 -2363
rect -515 -2369 -509 -2367
rect -505 -2363 -499 -2361
rect 547 -2362 553 -2360
rect 557 -2362 574 -2354
rect 578 -2356 595 -2354
rect 578 -2360 581 -2356
rect 585 -2360 595 -2356
rect 578 -2362 595 -2360
rect 613 -2356 619 -2354
rect 613 -2360 614 -2356
rect 618 -2360 619 -2356
rect 613 -2362 619 -2360
rect 623 -2356 629 -2354
rect 623 -2360 624 -2356
rect 628 -2360 629 -2356
rect 623 -2362 629 -2360
rect -505 -2367 -504 -2363
rect -500 -2367 -499 -2363
rect -505 -2369 -499 -2367
rect 35 -2536 41 -2534
rect 35 -2540 36 -2536
rect 40 -2540 41 -2536
rect 35 -2542 41 -2540
rect 45 -2536 62 -2534
rect 45 -2540 46 -2536
rect 50 -2540 62 -2536
rect 45 -2542 62 -2540
rect 66 -2536 83 -2534
rect 66 -2540 69 -2536
rect 73 -2540 83 -2536
rect 66 -2542 83 -2540
rect 87 -2536 104 -2534
rect 87 -2540 93 -2536
rect 97 -2540 104 -2536
rect 87 -2542 104 -2540
rect 108 -2542 146 -2534
rect 166 -2536 172 -2534
rect 166 -2540 167 -2536
rect 171 -2540 172 -2536
rect 166 -2542 172 -2540
rect 176 -2536 182 -2534
rect 176 -2540 177 -2536
rect 181 -2540 182 -2536
rect 176 -2542 182 -2540
rect 305 -2539 311 -2537
rect 305 -2543 306 -2539
rect 310 -2543 311 -2539
rect 305 -2545 311 -2543
rect 315 -2539 332 -2537
rect 315 -2543 316 -2539
rect 320 -2543 332 -2539
rect 315 -2545 332 -2543
rect 336 -2539 353 -2537
rect 336 -2543 339 -2539
rect 343 -2543 353 -2539
rect 336 -2545 353 -2543
rect 357 -2539 374 -2537
rect 357 -2543 363 -2539
rect 367 -2543 374 -2539
rect 357 -2545 374 -2543
rect 378 -2545 416 -2537
rect 436 -2539 442 -2537
rect 436 -2543 437 -2539
rect 441 -2543 442 -2539
rect 436 -2545 442 -2543
rect 446 -2539 452 -2537
rect 446 -2543 447 -2539
rect 451 -2543 452 -2539
rect 446 -2545 452 -2543
rect -580 -2647 -574 -2645
rect -580 -2651 -579 -2647
rect -575 -2651 -574 -2647
rect -580 -2653 -574 -2651
rect -570 -2653 -553 -2645
rect -549 -2647 -532 -2645
rect -549 -2651 -546 -2647
rect -542 -2651 -532 -2647
rect -549 -2653 -532 -2651
rect -514 -2647 -508 -2645
rect -514 -2651 -513 -2647
rect -509 -2651 -508 -2647
rect -514 -2653 -508 -2651
rect -504 -2647 -498 -2645
rect -504 -2651 -503 -2647
rect -499 -2651 -498 -2647
rect -504 -2653 -498 -2651
rect -583 -2739 -577 -2737
rect -583 -2743 -582 -2739
rect -578 -2743 -577 -2739
rect -583 -2745 -577 -2743
rect -573 -2745 -556 -2737
rect -552 -2739 -535 -2737
rect -552 -2743 -549 -2739
rect -545 -2743 -535 -2739
rect -552 -2745 -535 -2743
rect -517 -2739 -511 -2737
rect -517 -2743 -516 -2739
rect -512 -2743 -511 -2739
rect -517 -2745 -511 -2743
rect -507 -2739 -501 -2737
rect -507 -2743 -506 -2739
rect -502 -2743 -501 -2739
rect -507 -2745 -501 -2743
rect -82 -2806 -76 -2804
rect -82 -2810 -81 -2806
rect -77 -2810 -76 -2806
rect -82 -2812 -76 -2810
rect -72 -2812 -55 -2804
rect -51 -2806 -34 -2804
rect -51 -2810 -48 -2806
rect -44 -2810 -34 -2806
rect -51 -2812 -34 -2810
rect -16 -2806 -10 -2804
rect -16 -2810 -15 -2806
rect -11 -2810 -10 -2806
rect -16 -2812 -10 -2810
rect -6 -2806 0 -2804
rect -6 -2810 -5 -2806
rect -1 -2810 0 -2806
rect -6 -2812 0 -2810
rect -583 -2831 -577 -2829
rect -583 -2835 -582 -2831
rect -578 -2835 -577 -2831
rect -583 -2837 -577 -2835
rect -573 -2837 -556 -2829
rect -552 -2831 -535 -2829
rect -552 -2835 -549 -2831
rect -545 -2835 -535 -2831
rect -552 -2837 -535 -2835
rect -517 -2831 -511 -2829
rect -517 -2835 -516 -2831
rect -512 -2835 -511 -2831
rect -517 -2837 -511 -2835
rect -507 -2831 -501 -2829
rect -507 -2835 -506 -2831
rect -502 -2835 -501 -2831
rect -507 -2837 -501 -2835
rect -82 -2899 -76 -2897
rect -82 -2903 -81 -2899
rect -77 -2903 -76 -2899
rect -82 -2905 -76 -2903
rect -72 -2905 -55 -2897
rect -51 -2899 -34 -2897
rect -51 -2903 -48 -2899
rect -44 -2903 -34 -2899
rect -51 -2905 -34 -2903
rect -16 -2899 -10 -2897
rect -16 -2903 -15 -2899
rect -11 -2903 -10 -2899
rect -16 -2905 -10 -2903
rect -6 -2899 0 -2897
rect -6 -2903 -5 -2899
rect -1 -2903 0 -2899
rect -6 -2905 0 -2903
rect -583 -2923 -577 -2921
rect -583 -2927 -582 -2923
rect -578 -2927 -577 -2923
rect -583 -2929 -577 -2927
rect -573 -2929 -556 -2921
rect -552 -2923 -535 -2921
rect -552 -2927 -549 -2923
rect -545 -2927 -535 -2923
rect -552 -2929 -535 -2927
rect -517 -2923 -511 -2921
rect -517 -2927 -516 -2923
rect -512 -2927 -511 -2923
rect -517 -2929 -511 -2927
rect -507 -2923 -501 -2921
rect -507 -2927 -506 -2923
rect -502 -2927 -501 -2923
rect -507 -2929 -501 -2927
rect -82 -2991 -76 -2989
rect -82 -2995 -81 -2991
rect -77 -2995 -76 -2991
rect -82 -2997 -76 -2995
rect -72 -2997 -55 -2989
rect -51 -2991 -34 -2989
rect -51 -2995 -48 -2991
rect -44 -2995 -34 -2991
rect -51 -2997 -34 -2995
rect -16 -2991 -10 -2989
rect -16 -2995 -15 -2991
rect -11 -2995 -10 -2991
rect -16 -2997 -10 -2995
rect -6 -2991 0 -2989
rect -6 -2995 -5 -2991
rect -1 -2995 0 -2991
rect -6 -2997 0 -2995
rect -578 -3014 -572 -3012
rect -578 -3018 -577 -3014
rect -573 -3018 -572 -3014
rect -578 -3020 -572 -3018
rect -568 -3020 -551 -3012
rect -547 -3014 -530 -3012
rect -547 -3018 -544 -3014
rect -540 -3018 -530 -3014
rect -547 -3020 -530 -3018
rect -512 -3014 -506 -3012
rect -512 -3018 -511 -3014
rect -507 -3018 -506 -3014
rect -512 -3020 -506 -3018
rect -502 -3014 -496 -3012
rect -502 -3018 -501 -3014
rect -497 -3018 -496 -3014
rect -502 -3020 -496 -3018
rect -82 -3084 -76 -3082
rect -82 -3088 -81 -3084
rect -77 -3088 -76 -3084
rect -82 -3090 -76 -3088
rect -72 -3090 -55 -3082
rect -51 -3084 -34 -3082
rect -51 -3088 -48 -3084
rect -44 -3088 -34 -3084
rect -51 -3090 -34 -3088
rect -16 -3084 -10 -3082
rect -16 -3088 -15 -3084
rect -11 -3088 -10 -3084
rect -16 -3090 -10 -3088
rect -6 -3084 0 -3082
rect -6 -3088 -5 -3084
rect -1 -3088 0 -3084
rect -6 -3090 0 -3088
rect -581 -3106 -575 -3104
rect -581 -3110 -580 -3106
rect -576 -3110 -575 -3106
rect -581 -3112 -575 -3110
rect -571 -3112 -554 -3104
rect -550 -3106 -533 -3104
rect -550 -3110 -547 -3106
rect -543 -3110 -533 -3106
rect -550 -3112 -533 -3110
rect -515 -3106 -509 -3104
rect -515 -3110 -514 -3106
rect -510 -3110 -509 -3106
rect -515 -3112 -509 -3110
rect -505 -3106 -499 -3104
rect -505 -3110 -504 -3106
rect -500 -3110 -499 -3106
rect -505 -3112 -499 -3110
rect -581 -3198 -575 -3196
rect -581 -3202 -580 -3198
rect -576 -3202 -575 -3198
rect -581 -3204 -575 -3202
rect -571 -3204 -554 -3196
rect -550 -3198 -533 -3196
rect -550 -3202 -547 -3198
rect -543 -3202 -533 -3198
rect -550 -3204 -533 -3202
rect -515 -3198 -509 -3196
rect -515 -3202 -514 -3198
rect -510 -3202 -509 -3198
rect -515 -3204 -509 -3202
rect -505 -3198 -499 -3196
rect -505 -3202 -504 -3198
rect -500 -3202 -499 -3198
rect -505 -3204 -499 -3202
rect -581 -3290 -575 -3288
rect -581 -3294 -580 -3290
rect -576 -3294 -575 -3290
rect -581 -3296 -575 -3294
rect -571 -3296 -554 -3288
rect -550 -3290 -533 -3288
rect -550 -3294 -547 -3290
rect -543 -3294 -533 -3290
rect -550 -3296 -533 -3294
rect -515 -3290 -509 -3288
rect -515 -3294 -514 -3290
rect -510 -3294 -509 -3290
rect -515 -3296 -509 -3294
rect -505 -3290 -499 -3288
rect -505 -3294 -504 -3290
rect -500 -3294 -499 -3290
rect -505 -3296 -499 -3294
<< pdiffusion >>
rect -878 145 -872 147
rect -878 141 -877 145
rect -873 141 -872 145
rect -878 139 -872 141
rect -868 145 -862 147
rect -868 141 -867 145
rect -863 141 -862 145
rect -868 139 -862 141
rect -802 145 -796 147
rect -802 141 -801 145
rect -797 141 -796 145
rect -802 139 -796 141
rect -792 145 -775 147
rect -792 141 -791 145
rect -787 141 -775 145
rect -792 139 -775 141
rect -771 145 -754 147
rect -771 141 -768 145
rect -764 141 -754 145
rect -771 139 -754 141
rect -736 145 -730 147
rect -736 141 -735 145
rect -731 141 -730 145
rect -736 139 -730 141
rect -726 145 -720 147
rect -726 141 -725 145
rect -721 141 -720 145
rect -726 139 -720 141
rect -632 145 -626 147
rect -632 141 -631 145
rect -627 141 -626 145
rect -632 139 -626 141
rect -622 145 -605 147
rect -622 141 -621 145
rect -617 141 -605 145
rect -622 139 -605 141
rect -601 145 -584 147
rect -601 141 -598 145
rect -594 141 -584 145
rect -601 139 -584 141
rect -566 145 -560 147
rect -566 141 -565 145
rect -561 141 -560 145
rect -566 139 -560 141
rect -556 145 -550 147
rect -556 141 -555 145
rect -551 141 -550 145
rect -556 139 -550 141
rect -875 36 -869 38
rect -875 32 -874 36
rect -870 32 -869 36
rect -875 30 -869 32
rect -865 36 -859 38
rect -865 32 -864 36
rect -860 32 -859 36
rect -865 30 -859 32
rect -802 36 -796 38
rect -802 32 -801 36
rect -797 32 -796 36
rect -802 30 -796 32
rect -792 36 -775 38
rect -792 32 -791 36
rect -787 32 -775 36
rect -792 30 -775 32
rect -771 36 -754 38
rect -771 32 -768 36
rect -764 32 -754 36
rect -771 30 -754 32
rect -736 36 -730 38
rect -736 32 -735 36
rect -731 32 -730 36
rect -736 30 -730 32
rect -726 36 -720 38
rect -726 32 -725 36
rect -721 32 -720 36
rect -726 30 -720 32
rect -636 36 -630 38
rect -636 32 -635 36
rect -631 32 -630 36
rect -636 30 -630 32
rect -626 36 -609 38
rect -626 32 -625 36
rect -621 32 -609 36
rect -626 30 -609 32
rect -605 36 -588 38
rect -605 32 -602 36
rect -598 32 -588 36
rect -605 30 -588 32
rect -570 36 -564 38
rect -570 32 -569 36
rect -565 32 -564 36
rect -570 30 -564 32
rect -560 36 -554 38
rect -560 32 -559 36
rect -555 32 -554 36
rect -560 30 -554 32
rect -442 36 -436 38
rect -442 32 -441 36
rect -437 32 -436 36
rect -442 30 -436 32
rect -432 36 -426 38
rect -432 32 -431 36
rect -427 32 -426 36
rect -432 30 -426 32
rect -153 -18 -147 -16
rect -153 -22 -152 -18
rect -148 -22 -147 -18
rect -153 -24 -147 -22
rect -143 -18 -126 -16
rect -143 -22 -142 -18
rect -138 -22 -126 -18
rect -143 -24 -126 -22
rect -122 -18 -105 -16
rect -122 -22 -119 -18
rect -115 -22 -105 -18
rect -122 -24 -105 -22
rect 445 -18 451 -16
rect 445 -22 446 -18
rect 450 -22 451 -18
rect 445 -24 451 -22
rect 455 -18 472 -16
rect 455 -22 456 -18
rect 460 -22 472 -18
rect 455 -24 472 -22
rect 476 -18 493 -16
rect 476 -22 479 -18
rect 483 -22 493 -18
rect 476 -24 493 -22
rect 1324 -18 1330 -16
rect 1324 -22 1325 -18
rect 1329 -22 1330 -18
rect 1324 -24 1330 -22
rect 1334 -18 1351 -16
rect 1334 -22 1335 -18
rect 1339 -22 1351 -18
rect 1334 -24 1351 -22
rect 1355 -18 1372 -16
rect 1355 -22 1358 -18
rect 1362 -22 1372 -18
rect 1355 -24 1372 -22
rect 2092 -18 2098 -16
rect 2092 -22 2093 -18
rect 2097 -22 2098 -18
rect 2092 -24 2098 -22
rect 2102 -18 2119 -16
rect 2102 -22 2103 -18
rect 2107 -22 2119 -18
rect 2102 -24 2119 -22
rect 2123 -18 2140 -16
rect 2123 -22 2126 -18
rect 2130 -22 2140 -18
rect 2123 -24 2140 -22
rect -226 -66 -220 -64
rect -226 -70 -225 -66
rect -221 -70 -220 -66
rect -226 -72 -220 -70
rect -216 -66 -199 -64
rect -216 -70 -215 -66
rect -211 -70 -199 -66
rect -216 -72 -199 -70
rect -195 -66 -178 -64
rect -195 -70 -192 -66
rect -188 -70 -178 -66
rect 372 -66 378 -64
rect -195 -72 -178 -70
rect 372 -70 373 -66
rect 377 -70 378 -66
rect 372 -72 378 -70
rect 382 -66 399 -64
rect 382 -70 383 -66
rect 387 -70 399 -66
rect 382 -72 399 -70
rect 403 -66 420 -64
rect 403 -70 406 -66
rect 410 -70 420 -66
rect 1251 -66 1257 -64
rect 403 -72 420 -70
rect -52 -86 -46 -84
rect -52 -90 -51 -86
rect -47 -90 -46 -86
rect -52 -92 -46 -90
rect -42 -86 -25 -84
rect -42 -90 -41 -86
rect -37 -90 -25 -86
rect -42 -92 -25 -90
rect -21 -86 -4 -84
rect -21 -90 -18 -86
rect -14 -90 -4 -86
rect -21 -92 -4 -90
rect -580 -119 -574 -117
rect -580 -123 -579 -119
rect -575 -123 -574 -119
rect -580 -125 -574 -123
rect -570 -119 -553 -117
rect -570 -123 -569 -119
rect -565 -123 -553 -119
rect -570 -125 -553 -123
rect -549 -119 -532 -117
rect -549 -123 -546 -119
rect -542 -123 -532 -119
rect -549 -125 -532 -123
rect -514 -119 -508 -117
rect -514 -123 -513 -119
rect -509 -123 -508 -119
rect -514 -125 -508 -123
rect -504 -119 -498 -117
rect -504 -123 -503 -119
rect -499 -123 -498 -119
rect -504 -125 -498 -123
rect -138 -127 -132 -125
rect -138 -131 -137 -127
rect -133 -131 -132 -127
rect -138 -133 -132 -131
rect -128 -127 -111 -125
rect -128 -131 -127 -127
rect -123 -131 -111 -127
rect -128 -133 -111 -131
rect -107 -127 -90 -125
rect -107 -131 -104 -127
rect -100 -131 -90 -127
rect 1251 -70 1252 -66
rect 1256 -70 1257 -66
rect 1251 -72 1257 -70
rect 1261 -66 1278 -64
rect 1261 -70 1262 -66
rect 1266 -70 1278 -66
rect 1261 -72 1278 -70
rect 1282 -66 1299 -64
rect 1282 -70 1285 -66
rect 1289 -70 1299 -66
rect 2019 -66 2025 -64
rect 1282 -72 1299 -70
rect 546 -86 552 -84
rect 546 -90 547 -86
rect 551 -90 552 -86
rect 546 -92 552 -90
rect 556 -86 573 -84
rect 556 -90 557 -86
rect 561 -90 573 -86
rect 556 -92 573 -90
rect 577 -86 594 -84
rect 577 -90 580 -86
rect 584 -90 594 -86
rect 577 -92 594 -90
rect 460 -127 466 -125
rect -107 -133 -90 -131
rect 460 -131 461 -127
rect 465 -131 466 -127
rect 460 -133 466 -131
rect 470 -127 487 -125
rect 470 -131 471 -127
rect 475 -131 487 -127
rect 470 -133 487 -131
rect 491 -127 508 -125
rect 491 -131 494 -127
rect 498 -131 508 -127
rect 2019 -70 2020 -66
rect 2024 -70 2025 -66
rect 2019 -72 2025 -70
rect 2029 -66 2046 -64
rect 2029 -70 2030 -66
rect 2034 -70 2046 -66
rect 2029 -72 2046 -70
rect 2050 -66 2067 -64
rect 2050 -70 2053 -66
rect 2057 -70 2067 -66
rect 2050 -72 2067 -70
rect 1425 -86 1431 -84
rect 1425 -90 1426 -86
rect 1430 -90 1431 -86
rect 1425 -92 1431 -90
rect 1435 -86 1452 -84
rect 1435 -90 1436 -86
rect 1440 -90 1452 -86
rect 1435 -92 1452 -90
rect 1456 -86 1473 -84
rect 1456 -90 1459 -86
rect 1463 -90 1473 -86
rect 1456 -92 1473 -90
rect 1339 -127 1345 -125
rect 491 -133 508 -131
rect 1339 -131 1340 -127
rect 1344 -131 1345 -127
rect 1339 -133 1345 -131
rect 1349 -127 1366 -125
rect 1349 -131 1350 -127
rect 1354 -131 1366 -127
rect 1349 -133 1366 -131
rect 1370 -127 1387 -125
rect 1370 -131 1373 -127
rect 1377 -131 1387 -127
rect 2193 -86 2199 -84
rect 2193 -90 2194 -86
rect 2198 -90 2199 -86
rect 2193 -92 2199 -90
rect 2203 -86 2220 -84
rect 2203 -90 2204 -86
rect 2208 -90 2220 -86
rect 2203 -92 2220 -90
rect 2224 -86 2241 -84
rect 2224 -90 2227 -86
rect 2231 -90 2241 -86
rect 2224 -92 2241 -90
rect 2107 -127 2113 -125
rect 1370 -133 1387 -131
rect 2107 -131 2108 -127
rect 2112 -131 2113 -127
rect 2107 -133 2113 -131
rect 2117 -127 2134 -125
rect 2117 -131 2118 -127
rect 2122 -131 2134 -127
rect 2117 -133 2134 -131
rect 2138 -127 2155 -125
rect 2138 -131 2141 -127
rect 2145 -131 2155 -127
rect 2138 -133 2155 -131
rect -583 -211 -577 -209
rect -583 -215 -582 -211
rect -578 -215 -577 -211
rect -583 -217 -577 -215
rect -573 -211 -556 -209
rect -573 -215 -572 -211
rect -568 -215 -556 -211
rect -573 -217 -556 -215
rect -552 -211 -535 -209
rect -552 -215 -549 -211
rect -545 -215 -535 -211
rect -552 -217 -535 -215
rect -517 -211 -511 -209
rect -517 -215 -516 -211
rect -512 -215 -511 -211
rect -517 -217 -511 -215
rect -507 -211 -501 -209
rect -507 -215 -506 -211
rect -502 -215 -501 -211
rect -507 -217 -501 -215
rect -583 -303 -577 -301
rect -583 -307 -582 -303
rect -578 -307 -577 -303
rect -583 -309 -577 -307
rect -573 -303 -556 -301
rect -573 -307 -572 -303
rect -568 -307 -556 -303
rect -573 -309 -556 -307
rect -552 -303 -535 -301
rect -552 -307 -549 -303
rect -545 -307 -535 -303
rect -552 -309 -535 -307
rect -517 -303 -511 -301
rect -517 -307 -516 -303
rect -512 -307 -511 -303
rect -517 -309 -511 -307
rect -507 -303 -501 -301
rect -507 -307 -506 -303
rect -502 -307 -501 -303
rect -507 -309 -501 -307
rect 128 -321 134 -319
rect 128 -325 129 -321
rect 133 -325 134 -321
rect 128 -327 134 -325
rect 138 -321 155 -319
rect 138 -325 139 -321
rect 143 -325 155 -321
rect 138 -327 155 -325
rect 159 -321 176 -319
rect 159 -325 162 -321
rect 166 -325 176 -321
rect 159 -327 176 -325
rect 871 -324 877 -322
rect 871 -328 872 -324
rect 876 -328 877 -324
rect 871 -330 877 -328
rect 881 -324 898 -322
rect 881 -328 882 -324
rect 886 -328 898 -324
rect 881 -330 898 -328
rect 902 -324 919 -322
rect 902 -328 905 -324
rect 909 -328 919 -324
rect 902 -330 919 -328
rect 1630 -324 1636 -322
rect 1630 -328 1631 -324
rect 1635 -328 1636 -324
rect 1630 -330 1636 -328
rect 1640 -324 1657 -322
rect 1640 -328 1641 -324
rect 1645 -328 1657 -324
rect 1640 -330 1657 -328
rect 1661 -324 1678 -322
rect 1661 -328 1664 -324
rect 1668 -328 1678 -324
rect 1661 -330 1678 -328
rect 2366 -324 2372 -322
rect 2366 -328 2367 -324
rect 2371 -328 2372 -324
rect 2366 -330 2372 -328
rect 2376 -324 2393 -322
rect 2376 -328 2377 -324
rect 2381 -328 2393 -324
rect 2376 -330 2393 -328
rect 2397 -324 2414 -322
rect 2397 -328 2400 -324
rect 2404 -328 2414 -324
rect 2397 -330 2414 -328
rect -182 -369 -176 -367
rect -182 -373 -181 -369
rect -177 -373 -176 -369
rect -182 -375 -176 -373
rect -172 -369 -155 -367
rect -172 -373 -171 -369
rect -167 -373 -155 -369
rect -172 -375 -155 -373
rect -151 -369 -134 -367
rect -151 -373 -148 -369
rect -144 -373 -134 -369
rect -151 -375 -134 -373
rect 55 -369 61 -367
rect 55 -373 56 -369
rect 60 -373 61 -369
rect 55 -375 61 -373
rect 65 -369 82 -367
rect 65 -373 66 -369
rect 70 -373 82 -369
rect 65 -375 82 -373
rect 86 -369 103 -367
rect 86 -373 89 -369
rect 93 -373 103 -369
rect 561 -372 567 -370
rect 86 -375 103 -373
rect -583 -395 -577 -393
rect -583 -399 -582 -395
rect -578 -399 -577 -395
rect -583 -401 -577 -399
rect -573 -395 -556 -393
rect -573 -399 -572 -395
rect -568 -399 -556 -395
rect -573 -401 -556 -399
rect -552 -395 -535 -393
rect -552 -399 -549 -395
rect -545 -399 -535 -395
rect -552 -401 -535 -399
rect -517 -395 -511 -393
rect -517 -399 -516 -395
rect -512 -399 -511 -395
rect -517 -401 -511 -399
rect -507 -395 -501 -393
rect -507 -399 -506 -395
rect -502 -399 -501 -395
rect -507 -401 -501 -399
rect 561 -376 562 -372
rect 566 -376 567 -372
rect 561 -378 567 -376
rect 571 -372 588 -370
rect 571 -376 572 -372
rect 576 -376 588 -372
rect 571 -378 588 -376
rect 592 -372 609 -370
rect 592 -376 595 -372
rect 599 -376 609 -372
rect 592 -378 609 -376
rect 798 -372 804 -370
rect 798 -376 799 -372
rect 803 -376 804 -372
rect 798 -378 804 -376
rect 808 -372 825 -370
rect 808 -376 809 -372
rect 813 -376 825 -372
rect 808 -378 825 -376
rect 829 -372 846 -370
rect 829 -376 832 -372
rect 836 -376 846 -372
rect 1320 -372 1326 -370
rect 829 -378 846 -376
rect 229 -389 235 -387
rect 229 -393 230 -389
rect 234 -393 235 -389
rect 229 -395 235 -393
rect 239 -389 256 -387
rect 239 -393 240 -389
rect 244 -393 256 -389
rect 239 -395 256 -393
rect 260 -389 277 -387
rect 260 -393 263 -389
rect 267 -393 277 -389
rect 260 -395 277 -393
rect -255 -417 -249 -415
rect -255 -421 -254 -417
rect -250 -421 -249 -417
rect -255 -423 -249 -421
rect -245 -417 -228 -415
rect -245 -421 -244 -417
rect -240 -421 -228 -417
rect -245 -423 -228 -421
rect -224 -417 -207 -415
rect -224 -421 -221 -417
rect -217 -421 -207 -417
rect -224 -423 -207 -421
rect 143 -430 149 -428
rect 143 -434 144 -430
rect 148 -434 149 -430
rect -81 -437 -75 -435
rect -81 -441 -80 -437
rect -76 -441 -75 -437
rect -81 -443 -75 -441
rect -71 -437 -54 -435
rect -71 -441 -70 -437
rect -66 -441 -54 -437
rect -71 -443 -54 -441
rect -50 -437 -33 -435
rect 143 -436 149 -434
rect 153 -430 170 -428
rect 153 -434 154 -430
rect 158 -434 170 -430
rect 153 -436 170 -434
rect 174 -430 191 -428
rect 174 -434 177 -430
rect 181 -434 191 -430
rect 1320 -376 1321 -372
rect 1325 -376 1326 -372
rect 1320 -378 1326 -376
rect 1330 -372 1347 -370
rect 1330 -376 1331 -372
rect 1335 -376 1347 -372
rect 1330 -378 1347 -376
rect 1351 -372 1368 -370
rect 1351 -376 1354 -372
rect 1358 -376 1368 -372
rect 1351 -378 1368 -376
rect 1557 -372 1563 -370
rect 1557 -376 1558 -372
rect 1562 -376 1563 -372
rect 1557 -378 1563 -376
rect 1567 -372 1584 -370
rect 1567 -376 1568 -372
rect 1572 -376 1584 -372
rect 1567 -378 1584 -376
rect 1588 -372 1605 -370
rect 1588 -376 1591 -372
rect 1595 -376 1605 -372
rect 2056 -372 2062 -370
rect 1588 -378 1605 -376
rect 972 -392 978 -390
rect 972 -396 973 -392
rect 977 -396 978 -392
rect 972 -398 978 -396
rect 982 -392 999 -390
rect 982 -396 983 -392
rect 987 -396 999 -392
rect 982 -398 999 -396
rect 1003 -392 1020 -390
rect 1003 -396 1006 -392
rect 1010 -396 1020 -392
rect 1003 -398 1020 -396
rect 488 -420 494 -418
rect 488 -424 489 -420
rect 493 -424 494 -420
rect 488 -426 494 -424
rect 498 -420 515 -418
rect 498 -424 499 -420
rect 503 -424 515 -420
rect 498 -426 515 -424
rect 519 -420 536 -418
rect 519 -424 522 -420
rect 526 -424 536 -420
rect 519 -426 536 -424
rect 174 -436 191 -434
rect -50 -441 -47 -437
rect -43 -441 -33 -437
rect -50 -443 -33 -441
rect -167 -478 -161 -476
rect -167 -482 -166 -478
rect -162 -482 -161 -478
rect -167 -484 -161 -482
rect -157 -478 -140 -476
rect -157 -482 -156 -478
rect -152 -482 -140 -478
rect -157 -484 -140 -482
rect -136 -478 -119 -476
rect -136 -482 -133 -478
rect -129 -482 -119 -478
rect 886 -433 892 -431
rect 886 -437 887 -433
rect 891 -437 892 -433
rect 662 -440 668 -438
rect 662 -444 663 -440
rect 667 -444 668 -440
rect 662 -446 668 -444
rect 672 -440 689 -438
rect 672 -444 673 -440
rect 677 -444 689 -440
rect 672 -446 689 -444
rect 693 -440 710 -438
rect 886 -439 892 -437
rect 896 -433 913 -431
rect 896 -437 897 -433
rect 901 -437 913 -433
rect 896 -439 913 -437
rect 917 -433 934 -431
rect 917 -437 920 -433
rect 924 -437 934 -433
rect 2056 -376 2057 -372
rect 2061 -376 2062 -372
rect 2056 -378 2062 -376
rect 2066 -372 2083 -370
rect 2066 -376 2067 -372
rect 2071 -376 2083 -372
rect 2066 -378 2083 -376
rect 2087 -372 2104 -370
rect 2087 -376 2090 -372
rect 2094 -376 2104 -372
rect 2087 -378 2104 -376
rect 2293 -372 2299 -370
rect 2293 -376 2294 -372
rect 2298 -376 2299 -372
rect 2293 -378 2299 -376
rect 2303 -372 2320 -370
rect 2303 -376 2304 -372
rect 2308 -376 2320 -372
rect 2303 -378 2320 -376
rect 2324 -372 2341 -370
rect 2324 -376 2327 -372
rect 2331 -376 2341 -372
rect 2324 -378 2341 -376
rect 1731 -392 1737 -390
rect 1731 -396 1732 -392
rect 1736 -396 1737 -392
rect 1731 -398 1737 -396
rect 1741 -392 1758 -390
rect 1741 -396 1742 -392
rect 1746 -396 1758 -392
rect 1741 -398 1758 -396
rect 1762 -392 1779 -390
rect 1762 -396 1765 -392
rect 1769 -396 1779 -392
rect 1762 -398 1779 -396
rect 1247 -420 1253 -418
rect 1247 -424 1248 -420
rect 1252 -424 1253 -420
rect 1247 -426 1253 -424
rect 1257 -420 1274 -418
rect 1257 -424 1258 -420
rect 1262 -424 1274 -420
rect 1257 -426 1274 -424
rect 1278 -420 1295 -418
rect 1278 -424 1281 -420
rect 1285 -424 1295 -420
rect 1278 -426 1295 -424
rect 917 -439 934 -437
rect 693 -444 696 -440
rect 700 -444 710 -440
rect 693 -446 710 -444
rect -136 -484 -119 -482
rect -578 -486 -572 -484
rect -578 -490 -577 -486
rect -573 -490 -572 -486
rect -578 -492 -572 -490
rect -568 -486 -551 -484
rect -568 -490 -567 -486
rect -563 -490 -551 -486
rect -568 -492 -551 -490
rect -547 -486 -530 -484
rect -547 -490 -544 -486
rect -540 -490 -530 -486
rect -547 -492 -530 -490
rect -512 -486 -506 -484
rect -512 -490 -511 -486
rect -507 -490 -506 -486
rect -512 -492 -506 -490
rect -502 -486 -496 -484
rect -502 -490 -501 -486
rect -497 -490 -496 -486
rect -502 -492 -496 -490
rect 576 -481 582 -479
rect 576 -485 577 -481
rect 581 -485 582 -481
rect 576 -487 582 -485
rect 586 -481 603 -479
rect 586 -485 587 -481
rect 591 -485 603 -481
rect 586 -487 603 -485
rect 607 -481 624 -479
rect 607 -485 610 -481
rect 614 -485 624 -481
rect 1645 -433 1651 -431
rect 1645 -437 1646 -433
rect 1650 -437 1651 -433
rect 1421 -440 1427 -438
rect 1421 -444 1422 -440
rect 1426 -444 1427 -440
rect 1421 -446 1427 -444
rect 1431 -440 1448 -438
rect 1431 -444 1432 -440
rect 1436 -444 1448 -440
rect 1431 -446 1448 -444
rect 1452 -440 1469 -438
rect 1645 -439 1651 -437
rect 1655 -433 1672 -431
rect 1655 -437 1656 -433
rect 1660 -437 1672 -433
rect 1655 -439 1672 -437
rect 1676 -433 1693 -431
rect 1676 -437 1679 -433
rect 1683 -437 1693 -433
rect 2467 -392 2473 -390
rect 2467 -396 2468 -392
rect 2472 -396 2473 -392
rect 2467 -398 2473 -396
rect 2477 -392 2494 -390
rect 2477 -396 2478 -392
rect 2482 -396 2494 -392
rect 2477 -398 2494 -396
rect 2498 -392 2515 -390
rect 2498 -396 2501 -392
rect 2505 -396 2515 -392
rect 2498 -398 2515 -396
rect 1983 -420 1989 -418
rect 1983 -424 1984 -420
rect 1988 -424 1989 -420
rect 1983 -426 1989 -424
rect 1993 -420 2010 -418
rect 1993 -424 1994 -420
rect 1998 -424 2010 -420
rect 1993 -426 2010 -424
rect 2014 -420 2031 -418
rect 2014 -424 2017 -420
rect 2021 -424 2031 -420
rect 2014 -426 2031 -424
rect 1676 -439 1693 -437
rect 1452 -444 1455 -440
rect 1459 -444 1469 -440
rect 1452 -446 1469 -444
rect 607 -487 624 -485
rect 1335 -481 1341 -479
rect 1335 -485 1336 -481
rect 1340 -485 1341 -481
rect 1335 -487 1341 -485
rect 1345 -481 1362 -479
rect 1345 -485 1346 -481
rect 1350 -485 1362 -481
rect 1345 -487 1362 -485
rect 1366 -481 1383 -479
rect 1366 -485 1369 -481
rect 1373 -485 1383 -481
rect 2381 -433 2387 -431
rect 2381 -437 2382 -433
rect 2386 -437 2387 -433
rect 2157 -440 2163 -438
rect 2157 -444 2158 -440
rect 2162 -444 2163 -440
rect 2157 -446 2163 -444
rect 2167 -440 2184 -438
rect 2167 -444 2168 -440
rect 2172 -444 2184 -440
rect 2167 -446 2184 -444
rect 2188 -440 2205 -438
rect 2381 -439 2387 -437
rect 2391 -433 2408 -431
rect 2391 -437 2392 -433
rect 2396 -437 2408 -433
rect 2391 -439 2408 -437
rect 2412 -433 2429 -431
rect 2412 -437 2415 -433
rect 2419 -437 2429 -433
rect 2412 -439 2429 -437
rect 2188 -444 2191 -440
rect 2195 -444 2205 -440
rect 2188 -446 2205 -444
rect 1366 -487 1383 -485
rect 2071 -481 2077 -479
rect 2071 -485 2072 -481
rect 2076 -485 2077 -481
rect 2071 -487 2077 -485
rect 2081 -481 2098 -479
rect 2081 -485 2082 -481
rect 2086 -485 2098 -481
rect 2081 -487 2098 -485
rect 2102 -481 2119 -479
rect 2102 -485 2105 -481
rect 2109 -485 2119 -481
rect 2102 -487 2119 -485
rect 115 -536 121 -534
rect 115 -540 116 -536
rect 120 -540 121 -536
rect 115 -542 121 -540
rect 125 -536 142 -534
rect 125 -540 126 -536
rect 130 -540 142 -536
rect 125 -542 142 -540
rect 146 -536 163 -534
rect 146 -540 149 -536
rect 153 -540 163 -536
rect 146 -542 163 -540
rect 181 -536 187 -534
rect 181 -540 182 -536
rect 186 -540 187 -536
rect 181 -542 187 -540
rect 191 -536 197 -534
rect 191 -540 192 -536
rect 196 -540 197 -536
rect 191 -542 197 -540
rect 274 -536 280 -534
rect 274 -540 275 -536
rect 279 -540 280 -536
rect 274 -542 280 -540
rect 284 -542 301 -534
rect 305 -536 322 -534
rect 305 -540 310 -536
rect 314 -540 322 -536
rect 305 -542 322 -540
rect 342 -536 348 -534
rect 342 -540 343 -536
rect 347 -540 348 -536
rect 342 -542 348 -540
rect 352 -536 358 -534
rect 352 -540 353 -536
rect 357 -540 358 -536
rect 858 -539 864 -537
rect 352 -542 358 -540
rect -581 -578 -575 -576
rect -581 -582 -580 -578
rect -576 -582 -575 -578
rect -581 -584 -575 -582
rect -571 -578 -554 -576
rect -571 -582 -570 -578
rect -566 -582 -554 -578
rect -571 -584 -554 -582
rect -550 -578 -533 -576
rect -550 -582 -547 -578
rect -543 -582 -533 -578
rect -550 -584 -533 -582
rect -515 -578 -509 -576
rect -515 -582 -514 -578
rect -510 -582 -509 -578
rect -515 -584 -509 -582
rect -505 -578 -499 -576
rect -505 -582 -504 -578
rect -500 -582 -499 -578
rect -505 -584 -499 -582
rect -196 -587 -190 -585
rect -196 -591 -195 -587
rect -191 -591 -190 -587
rect -196 -593 -190 -591
rect -186 -587 -169 -585
rect -186 -591 -185 -587
rect -181 -591 -169 -587
rect -186 -593 -169 -591
rect -165 -587 -148 -585
rect -165 -591 -162 -587
rect -158 -591 -148 -587
rect -165 -593 -148 -591
rect -130 -587 -124 -585
rect -130 -591 -129 -587
rect -125 -591 -124 -587
rect -130 -593 -124 -591
rect -120 -587 -114 -585
rect 858 -543 859 -539
rect 863 -543 864 -539
rect 858 -545 864 -543
rect 868 -539 885 -537
rect 868 -543 869 -539
rect 873 -543 885 -539
rect 868 -545 885 -543
rect 889 -539 906 -537
rect 889 -543 892 -539
rect 896 -543 906 -539
rect 889 -545 906 -543
rect 924 -539 930 -537
rect 924 -543 925 -539
rect 929 -543 930 -539
rect 924 -545 930 -543
rect 934 -539 940 -537
rect 934 -543 935 -539
rect 939 -543 940 -539
rect 934 -545 940 -543
rect 1017 -539 1023 -537
rect 1017 -543 1018 -539
rect 1022 -543 1023 -539
rect 1017 -545 1023 -543
rect 1027 -545 1044 -537
rect 1048 -539 1065 -537
rect 1048 -543 1053 -539
rect 1057 -543 1065 -539
rect 1048 -545 1065 -543
rect 1085 -539 1091 -537
rect 1085 -543 1086 -539
rect 1090 -543 1091 -539
rect 1085 -545 1091 -543
rect 1095 -539 1101 -537
rect 1095 -543 1096 -539
rect 1100 -543 1101 -539
rect 1617 -539 1623 -537
rect 1095 -545 1101 -543
rect 1617 -543 1618 -539
rect 1622 -543 1623 -539
rect 1617 -545 1623 -543
rect 1627 -539 1644 -537
rect 1627 -543 1628 -539
rect 1632 -543 1644 -539
rect 1627 -545 1644 -543
rect 1648 -539 1665 -537
rect 1648 -543 1651 -539
rect 1655 -543 1665 -539
rect 1648 -545 1665 -543
rect 1683 -539 1689 -537
rect 1683 -543 1684 -539
rect 1688 -543 1689 -539
rect 1683 -545 1689 -543
rect 1693 -539 1699 -537
rect 1693 -543 1694 -539
rect 1698 -543 1699 -539
rect 1693 -545 1699 -543
rect 1776 -539 1782 -537
rect 1776 -543 1777 -539
rect 1781 -543 1782 -539
rect 1776 -545 1782 -543
rect 1786 -545 1803 -537
rect 1807 -539 1824 -537
rect 1807 -543 1812 -539
rect 1816 -543 1824 -539
rect 1807 -545 1824 -543
rect 1844 -539 1850 -537
rect 1844 -543 1845 -539
rect 1849 -543 1850 -539
rect 1844 -545 1850 -543
rect 1854 -539 1860 -537
rect 1854 -543 1855 -539
rect 1859 -543 1860 -539
rect 2353 -539 2359 -537
rect 1854 -545 1860 -543
rect 2353 -543 2354 -539
rect 2358 -543 2359 -539
rect 2353 -545 2359 -543
rect 2363 -539 2380 -537
rect 2363 -543 2364 -539
rect 2368 -543 2380 -539
rect 2363 -545 2380 -543
rect 2384 -539 2401 -537
rect 2384 -543 2387 -539
rect 2391 -543 2401 -539
rect 2384 -545 2401 -543
rect 2419 -539 2425 -537
rect 2419 -543 2420 -539
rect 2424 -543 2425 -539
rect 2419 -545 2425 -543
rect 2429 -539 2435 -537
rect 2429 -543 2430 -539
rect 2434 -543 2435 -539
rect 2429 -545 2435 -543
rect 2512 -539 2518 -537
rect 2512 -543 2513 -539
rect 2517 -543 2518 -539
rect 2512 -545 2518 -543
rect 2522 -545 2539 -537
rect 2543 -539 2560 -537
rect 2543 -543 2548 -539
rect 2552 -543 2560 -539
rect 2543 -545 2560 -543
rect 2580 -539 2586 -537
rect 2580 -543 2581 -539
rect 2585 -543 2586 -539
rect 2580 -545 2586 -543
rect 2590 -539 2596 -537
rect 2590 -543 2591 -539
rect 2595 -543 2596 -539
rect 2590 -545 2596 -543
rect -120 -591 -119 -587
rect -115 -591 -114 -587
rect 547 -590 553 -588
rect -120 -593 -114 -591
rect 547 -594 548 -590
rect 552 -594 553 -590
rect 547 -596 553 -594
rect 557 -590 574 -588
rect 557 -594 558 -590
rect 562 -594 574 -590
rect 557 -596 574 -594
rect 578 -590 595 -588
rect 578 -594 581 -590
rect 585 -594 595 -590
rect 578 -596 595 -594
rect 613 -590 619 -588
rect 613 -594 614 -590
rect 618 -594 619 -590
rect 613 -596 619 -594
rect 623 -590 629 -588
rect 623 -594 624 -590
rect 628 -594 629 -590
rect 1306 -590 1312 -588
rect 623 -596 629 -594
rect 1306 -594 1307 -590
rect 1311 -594 1312 -590
rect 1306 -596 1312 -594
rect 1316 -590 1333 -588
rect 1316 -594 1317 -590
rect 1321 -594 1333 -590
rect 1316 -596 1333 -594
rect 1337 -590 1354 -588
rect 1337 -594 1340 -590
rect 1344 -594 1354 -590
rect 1337 -596 1354 -594
rect 1372 -590 1378 -588
rect 1372 -594 1373 -590
rect 1377 -594 1378 -590
rect 1372 -596 1378 -594
rect 1382 -590 1388 -588
rect 1382 -594 1383 -590
rect 1387 -594 1388 -590
rect 2042 -590 2048 -588
rect 1382 -596 1388 -594
rect 2042 -594 2043 -590
rect 2047 -594 2048 -590
rect 2042 -596 2048 -594
rect 2052 -590 2069 -588
rect 2052 -594 2053 -590
rect 2057 -594 2069 -590
rect 2052 -596 2069 -594
rect 2073 -590 2090 -588
rect 2073 -594 2076 -590
rect 2080 -594 2090 -590
rect 2073 -596 2090 -594
rect 2108 -590 2114 -588
rect 2108 -594 2109 -590
rect 2113 -594 2114 -590
rect 2108 -596 2114 -594
rect 2118 -590 2124 -588
rect 2118 -594 2119 -590
rect 2123 -594 2124 -590
rect 2118 -596 2124 -594
rect -581 -670 -575 -668
rect -581 -674 -580 -670
rect -576 -674 -575 -670
rect -581 -676 -575 -674
rect -571 -670 -554 -668
rect -571 -674 -570 -670
rect -566 -674 -554 -670
rect -571 -676 -554 -674
rect -550 -670 -533 -668
rect -550 -674 -547 -670
rect -543 -674 -533 -670
rect -550 -676 -533 -674
rect -515 -670 -509 -668
rect -515 -674 -514 -670
rect -510 -674 -509 -670
rect -515 -676 -509 -674
rect -505 -670 -499 -668
rect -505 -674 -504 -670
rect -500 -674 -499 -670
rect -505 -676 -499 -674
rect -581 -762 -575 -760
rect -581 -766 -580 -762
rect -576 -766 -575 -762
rect -581 -768 -575 -766
rect -571 -762 -554 -760
rect -571 -766 -570 -762
rect -566 -766 -554 -762
rect -571 -768 -554 -766
rect -550 -762 -533 -760
rect -550 -766 -547 -762
rect -543 -766 -533 -762
rect -550 -768 -533 -766
rect -515 -762 -509 -760
rect -515 -766 -514 -762
rect -510 -766 -509 -762
rect -515 -768 -509 -766
rect -505 -762 -499 -760
rect -505 -766 -504 -762
rect -500 -766 -499 -762
rect -505 -768 -499 -766
rect -124 -811 -118 -809
rect -124 -815 -123 -811
rect -119 -815 -118 -811
rect -124 -817 -118 -815
rect -114 -811 -97 -809
rect -114 -815 -113 -811
rect -109 -815 -97 -811
rect -114 -817 -97 -815
rect -93 -811 -76 -809
rect -93 -815 -90 -811
rect -86 -815 -76 -811
rect -93 -817 -76 -815
rect 474 -811 480 -809
rect 474 -815 475 -811
rect 479 -815 480 -811
rect 474 -817 480 -815
rect 484 -811 501 -809
rect 484 -815 485 -811
rect 489 -815 501 -811
rect 484 -817 501 -815
rect 505 -811 522 -809
rect 505 -815 508 -811
rect 512 -815 522 -811
rect 505 -817 522 -815
rect 1353 -811 1359 -809
rect 1353 -815 1354 -811
rect 1358 -815 1359 -811
rect 1353 -817 1359 -815
rect 1363 -811 1380 -809
rect 1363 -815 1364 -811
rect 1368 -815 1380 -811
rect 1363 -817 1380 -815
rect 1384 -811 1401 -809
rect 1384 -815 1387 -811
rect 1391 -815 1401 -811
rect 1384 -817 1401 -815
rect 2121 -811 2127 -809
rect 2121 -815 2122 -811
rect 2126 -815 2127 -811
rect 2121 -817 2127 -815
rect 2131 -811 2148 -809
rect 2131 -815 2132 -811
rect 2136 -815 2148 -811
rect 2131 -817 2148 -815
rect 2152 -811 2169 -809
rect 2152 -815 2155 -811
rect 2159 -815 2169 -811
rect 2152 -817 2169 -815
rect -197 -859 -191 -857
rect -197 -863 -196 -859
rect -192 -863 -191 -859
rect -197 -865 -191 -863
rect -187 -859 -170 -857
rect -187 -863 -186 -859
rect -182 -863 -170 -859
rect -187 -865 -170 -863
rect -166 -859 -149 -857
rect -166 -863 -163 -859
rect -159 -863 -149 -859
rect 401 -859 407 -857
rect -166 -865 -149 -863
rect 401 -863 402 -859
rect 406 -863 407 -859
rect 401 -865 407 -863
rect 411 -859 428 -857
rect 411 -863 412 -859
rect 416 -863 428 -859
rect 411 -865 428 -863
rect 432 -859 449 -857
rect 432 -863 435 -859
rect 439 -863 449 -859
rect 1280 -859 1286 -857
rect 432 -865 449 -863
rect -23 -879 -17 -877
rect -23 -883 -22 -879
rect -18 -883 -17 -879
rect -23 -885 -17 -883
rect -13 -879 4 -877
rect -13 -883 -12 -879
rect -8 -883 4 -879
rect -13 -885 4 -883
rect 8 -879 25 -877
rect 8 -883 11 -879
rect 15 -883 25 -879
rect 8 -885 25 -883
rect -580 -912 -574 -910
rect -580 -916 -579 -912
rect -575 -916 -574 -912
rect -580 -918 -574 -916
rect -570 -912 -553 -910
rect -570 -916 -569 -912
rect -565 -916 -553 -912
rect -570 -918 -553 -916
rect -549 -912 -532 -910
rect -549 -916 -546 -912
rect -542 -916 -532 -912
rect -549 -918 -532 -916
rect -514 -912 -508 -910
rect -514 -916 -513 -912
rect -509 -916 -508 -912
rect -514 -918 -508 -916
rect -504 -912 -498 -910
rect -504 -916 -503 -912
rect -499 -916 -498 -912
rect -504 -918 -498 -916
rect -109 -920 -103 -918
rect -109 -924 -108 -920
rect -104 -924 -103 -920
rect -109 -926 -103 -924
rect -99 -920 -82 -918
rect -99 -924 -98 -920
rect -94 -924 -82 -920
rect -99 -926 -82 -924
rect -78 -920 -61 -918
rect -78 -924 -75 -920
rect -71 -924 -61 -920
rect 1280 -863 1281 -859
rect 1285 -863 1286 -859
rect 1280 -865 1286 -863
rect 1290 -859 1307 -857
rect 1290 -863 1291 -859
rect 1295 -863 1307 -859
rect 1290 -865 1307 -863
rect 1311 -859 1328 -857
rect 1311 -863 1314 -859
rect 1318 -863 1328 -859
rect 2048 -859 2054 -857
rect 1311 -865 1328 -863
rect 575 -879 581 -877
rect 575 -883 576 -879
rect 580 -883 581 -879
rect 575 -885 581 -883
rect 585 -879 602 -877
rect 585 -883 586 -879
rect 590 -883 602 -879
rect 585 -885 602 -883
rect 606 -879 623 -877
rect 606 -883 609 -879
rect 613 -883 623 -879
rect 606 -885 623 -883
rect 489 -920 495 -918
rect -78 -926 -61 -924
rect 489 -924 490 -920
rect 494 -924 495 -920
rect 489 -926 495 -924
rect 499 -920 516 -918
rect 499 -924 500 -920
rect 504 -924 516 -920
rect 499 -926 516 -924
rect 520 -920 537 -918
rect 520 -924 523 -920
rect 527 -924 537 -920
rect 2048 -863 2049 -859
rect 2053 -863 2054 -859
rect 2048 -865 2054 -863
rect 2058 -859 2075 -857
rect 2058 -863 2059 -859
rect 2063 -863 2075 -859
rect 2058 -865 2075 -863
rect 2079 -859 2096 -857
rect 2079 -863 2082 -859
rect 2086 -863 2096 -859
rect 2079 -865 2096 -863
rect 1454 -879 1460 -877
rect 1454 -883 1455 -879
rect 1459 -883 1460 -879
rect 1454 -885 1460 -883
rect 1464 -879 1481 -877
rect 1464 -883 1465 -879
rect 1469 -883 1481 -879
rect 1464 -885 1481 -883
rect 1485 -879 1502 -877
rect 1485 -883 1488 -879
rect 1492 -883 1502 -879
rect 1485 -885 1502 -883
rect 1368 -920 1374 -918
rect 520 -926 537 -924
rect 1368 -924 1369 -920
rect 1373 -924 1374 -920
rect 1368 -926 1374 -924
rect 1378 -920 1395 -918
rect 1378 -924 1379 -920
rect 1383 -924 1395 -920
rect 1378 -926 1395 -924
rect 1399 -920 1416 -918
rect 1399 -924 1402 -920
rect 1406 -924 1416 -920
rect 2222 -879 2228 -877
rect 2222 -883 2223 -879
rect 2227 -883 2228 -879
rect 2222 -885 2228 -883
rect 2232 -879 2249 -877
rect 2232 -883 2233 -879
rect 2237 -883 2249 -879
rect 2232 -885 2249 -883
rect 2253 -879 2270 -877
rect 2253 -883 2256 -879
rect 2260 -883 2270 -879
rect 2253 -885 2270 -883
rect 2136 -920 2142 -918
rect 1399 -926 1416 -924
rect 2136 -924 2137 -920
rect 2141 -924 2142 -920
rect 2136 -926 2142 -924
rect 2146 -920 2163 -918
rect 2146 -924 2147 -920
rect 2151 -924 2163 -920
rect 2146 -926 2163 -924
rect 2167 -920 2184 -918
rect 2167 -924 2170 -920
rect 2174 -924 2184 -920
rect 2167 -926 2184 -924
rect -583 -1004 -577 -1002
rect -583 -1008 -582 -1004
rect -578 -1008 -577 -1004
rect -583 -1010 -577 -1008
rect -573 -1004 -556 -1002
rect -573 -1008 -572 -1004
rect -568 -1008 -556 -1004
rect -573 -1010 -556 -1008
rect -552 -1004 -535 -1002
rect -552 -1008 -549 -1004
rect -545 -1008 -535 -1004
rect -552 -1010 -535 -1008
rect -517 -1004 -511 -1002
rect -517 -1008 -516 -1004
rect -512 -1008 -511 -1004
rect -517 -1010 -511 -1008
rect -507 -1004 -501 -1002
rect -507 -1008 -506 -1004
rect -502 -1008 -501 -1004
rect -507 -1010 -501 -1008
rect -583 -1096 -577 -1094
rect -583 -1100 -582 -1096
rect -578 -1100 -577 -1096
rect -583 -1102 -577 -1100
rect -573 -1096 -556 -1094
rect -573 -1100 -572 -1096
rect -568 -1100 -556 -1096
rect -573 -1102 -556 -1100
rect -552 -1096 -535 -1094
rect -552 -1100 -549 -1096
rect -545 -1100 -535 -1096
rect -552 -1102 -535 -1100
rect -517 -1096 -511 -1094
rect -517 -1100 -516 -1096
rect -512 -1100 -511 -1096
rect -517 -1102 -511 -1100
rect -507 -1096 -501 -1094
rect -507 -1100 -506 -1096
rect -502 -1100 -501 -1096
rect -507 -1102 -501 -1100
rect 157 -1114 163 -1112
rect 157 -1118 158 -1114
rect 162 -1118 163 -1114
rect 157 -1120 163 -1118
rect 167 -1114 184 -1112
rect 167 -1118 168 -1114
rect 172 -1118 184 -1114
rect 167 -1120 184 -1118
rect 188 -1114 205 -1112
rect 188 -1118 191 -1114
rect 195 -1118 205 -1114
rect 188 -1120 205 -1118
rect 900 -1117 906 -1115
rect 900 -1121 901 -1117
rect 905 -1121 906 -1117
rect 900 -1123 906 -1121
rect 910 -1117 927 -1115
rect 910 -1121 911 -1117
rect 915 -1121 927 -1117
rect 910 -1123 927 -1121
rect 931 -1117 948 -1115
rect 931 -1121 934 -1117
rect 938 -1121 948 -1117
rect 931 -1123 948 -1121
rect 1659 -1117 1665 -1115
rect 1659 -1121 1660 -1117
rect 1664 -1121 1665 -1117
rect 1659 -1123 1665 -1121
rect 1669 -1117 1686 -1115
rect 1669 -1121 1670 -1117
rect 1674 -1121 1686 -1117
rect 1669 -1123 1686 -1121
rect 1690 -1117 1707 -1115
rect 1690 -1121 1693 -1117
rect 1697 -1121 1707 -1117
rect 1690 -1123 1707 -1121
rect 2395 -1117 2401 -1115
rect 2395 -1121 2396 -1117
rect 2400 -1121 2401 -1117
rect 2395 -1123 2401 -1121
rect 2405 -1117 2422 -1115
rect 2405 -1121 2406 -1117
rect 2410 -1121 2422 -1117
rect 2405 -1123 2422 -1121
rect 2426 -1117 2443 -1115
rect 2426 -1121 2429 -1117
rect 2433 -1121 2443 -1117
rect 2426 -1123 2443 -1121
rect -153 -1162 -147 -1160
rect -153 -1166 -152 -1162
rect -148 -1166 -147 -1162
rect -153 -1168 -147 -1166
rect -143 -1162 -126 -1160
rect -143 -1166 -142 -1162
rect -138 -1166 -126 -1162
rect -143 -1168 -126 -1166
rect -122 -1162 -105 -1160
rect -122 -1166 -119 -1162
rect -115 -1166 -105 -1162
rect -122 -1168 -105 -1166
rect 84 -1162 90 -1160
rect 84 -1166 85 -1162
rect 89 -1166 90 -1162
rect 84 -1168 90 -1166
rect 94 -1162 111 -1160
rect 94 -1166 95 -1162
rect 99 -1166 111 -1162
rect 94 -1168 111 -1166
rect 115 -1162 132 -1160
rect 115 -1166 118 -1162
rect 122 -1166 132 -1162
rect 590 -1165 596 -1163
rect 115 -1168 132 -1166
rect -583 -1188 -577 -1186
rect -583 -1192 -582 -1188
rect -578 -1192 -577 -1188
rect -583 -1194 -577 -1192
rect -573 -1188 -556 -1186
rect -573 -1192 -572 -1188
rect -568 -1192 -556 -1188
rect -573 -1194 -556 -1192
rect -552 -1188 -535 -1186
rect -552 -1192 -549 -1188
rect -545 -1192 -535 -1188
rect -552 -1194 -535 -1192
rect -517 -1188 -511 -1186
rect -517 -1192 -516 -1188
rect -512 -1192 -511 -1188
rect -517 -1194 -511 -1192
rect -507 -1188 -501 -1186
rect -507 -1192 -506 -1188
rect -502 -1192 -501 -1188
rect -507 -1194 -501 -1192
rect 590 -1169 591 -1165
rect 595 -1169 596 -1165
rect 590 -1171 596 -1169
rect 600 -1165 617 -1163
rect 600 -1169 601 -1165
rect 605 -1169 617 -1165
rect 600 -1171 617 -1169
rect 621 -1165 638 -1163
rect 621 -1169 624 -1165
rect 628 -1169 638 -1165
rect 621 -1171 638 -1169
rect 827 -1165 833 -1163
rect 827 -1169 828 -1165
rect 832 -1169 833 -1165
rect 827 -1171 833 -1169
rect 837 -1165 854 -1163
rect 837 -1169 838 -1165
rect 842 -1169 854 -1165
rect 837 -1171 854 -1169
rect 858 -1165 875 -1163
rect 858 -1169 861 -1165
rect 865 -1169 875 -1165
rect 1349 -1165 1355 -1163
rect 858 -1171 875 -1169
rect 258 -1182 264 -1180
rect 258 -1186 259 -1182
rect 263 -1186 264 -1182
rect 258 -1188 264 -1186
rect 268 -1182 285 -1180
rect 268 -1186 269 -1182
rect 273 -1186 285 -1182
rect 268 -1188 285 -1186
rect 289 -1182 306 -1180
rect 289 -1186 292 -1182
rect 296 -1186 306 -1182
rect 289 -1188 306 -1186
rect -226 -1210 -220 -1208
rect -226 -1214 -225 -1210
rect -221 -1214 -220 -1210
rect -226 -1216 -220 -1214
rect -216 -1210 -199 -1208
rect -216 -1214 -215 -1210
rect -211 -1214 -199 -1210
rect -216 -1216 -199 -1214
rect -195 -1210 -178 -1208
rect -195 -1214 -192 -1210
rect -188 -1214 -178 -1210
rect -195 -1216 -178 -1214
rect 172 -1223 178 -1221
rect 172 -1227 173 -1223
rect 177 -1227 178 -1223
rect -52 -1230 -46 -1228
rect -52 -1234 -51 -1230
rect -47 -1234 -46 -1230
rect -52 -1236 -46 -1234
rect -42 -1230 -25 -1228
rect -42 -1234 -41 -1230
rect -37 -1234 -25 -1230
rect -42 -1236 -25 -1234
rect -21 -1230 -4 -1228
rect 172 -1229 178 -1227
rect 182 -1223 199 -1221
rect 182 -1227 183 -1223
rect 187 -1227 199 -1223
rect 182 -1229 199 -1227
rect 203 -1223 220 -1221
rect 203 -1227 206 -1223
rect 210 -1227 220 -1223
rect 1349 -1169 1350 -1165
rect 1354 -1169 1355 -1165
rect 1349 -1171 1355 -1169
rect 1359 -1165 1376 -1163
rect 1359 -1169 1360 -1165
rect 1364 -1169 1376 -1165
rect 1359 -1171 1376 -1169
rect 1380 -1165 1397 -1163
rect 1380 -1169 1383 -1165
rect 1387 -1169 1397 -1165
rect 1380 -1171 1397 -1169
rect 1586 -1165 1592 -1163
rect 1586 -1169 1587 -1165
rect 1591 -1169 1592 -1165
rect 1586 -1171 1592 -1169
rect 1596 -1165 1613 -1163
rect 1596 -1169 1597 -1165
rect 1601 -1169 1613 -1165
rect 1596 -1171 1613 -1169
rect 1617 -1165 1634 -1163
rect 1617 -1169 1620 -1165
rect 1624 -1169 1634 -1165
rect 2085 -1165 2091 -1163
rect 1617 -1171 1634 -1169
rect 1001 -1185 1007 -1183
rect 1001 -1189 1002 -1185
rect 1006 -1189 1007 -1185
rect 1001 -1191 1007 -1189
rect 1011 -1185 1028 -1183
rect 1011 -1189 1012 -1185
rect 1016 -1189 1028 -1185
rect 1011 -1191 1028 -1189
rect 1032 -1185 1049 -1183
rect 1032 -1189 1035 -1185
rect 1039 -1189 1049 -1185
rect 1032 -1191 1049 -1189
rect 517 -1213 523 -1211
rect 517 -1217 518 -1213
rect 522 -1217 523 -1213
rect 517 -1219 523 -1217
rect 527 -1213 544 -1211
rect 527 -1217 528 -1213
rect 532 -1217 544 -1213
rect 527 -1219 544 -1217
rect 548 -1213 565 -1211
rect 548 -1217 551 -1213
rect 555 -1217 565 -1213
rect 548 -1219 565 -1217
rect 203 -1229 220 -1227
rect -21 -1234 -18 -1230
rect -14 -1234 -4 -1230
rect -21 -1236 -4 -1234
rect -138 -1271 -132 -1269
rect -138 -1275 -137 -1271
rect -133 -1275 -132 -1271
rect -138 -1277 -132 -1275
rect -128 -1271 -111 -1269
rect -128 -1275 -127 -1271
rect -123 -1275 -111 -1271
rect -128 -1277 -111 -1275
rect -107 -1271 -90 -1269
rect -107 -1275 -104 -1271
rect -100 -1275 -90 -1271
rect 915 -1226 921 -1224
rect 915 -1230 916 -1226
rect 920 -1230 921 -1226
rect 691 -1233 697 -1231
rect 691 -1237 692 -1233
rect 696 -1237 697 -1233
rect 691 -1239 697 -1237
rect 701 -1233 718 -1231
rect 701 -1237 702 -1233
rect 706 -1237 718 -1233
rect 701 -1239 718 -1237
rect 722 -1233 739 -1231
rect 915 -1232 921 -1230
rect 925 -1226 942 -1224
rect 925 -1230 926 -1226
rect 930 -1230 942 -1226
rect 925 -1232 942 -1230
rect 946 -1226 963 -1224
rect 946 -1230 949 -1226
rect 953 -1230 963 -1226
rect 2085 -1169 2086 -1165
rect 2090 -1169 2091 -1165
rect 2085 -1171 2091 -1169
rect 2095 -1165 2112 -1163
rect 2095 -1169 2096 -1165
rect 2100 -1169 2112 -1165
rect 2095 -1171 2112 -1169
rect 2116 -1165 2133 -1163
rect 2116 -1169 2119 -1165
rect 2123 -1169 2133 -1165
rect 2116 -1171 2133 -1169
rect 2322 -1165 2328 -1163
rect 2322 -1169 2323 -1165
rect 2327 -1169 2328 -1165
rect 2322 -1171 2328 -1169
rect 2332 -1165 2349 -1163
rect 2332 -1169 2333 -1165
rect 2337 -1169 2349 -1165
rect 2332 -1171 2349 -1169
rect 2353 -1165 2370 -1163
rect 2353 -1169 2356 -1165
rect 2360 -1169 2370 -1165
rect 2353 -1171 2370 -1169
rect 1760 -1185 1766 -1183
rect 1760 -1189 1761 -1185
rect 1765 -1189 1766 -1185
rect 1760 -1191 1766 -1189
rect 1770 -1185 1787 -1183
rect 1770 -1189 1771 -1185
rect 1775 -1189 1787 -1185
rect 1770 -1191 1787 -1189
rect 1791 -1185 1808 -1183
rect 1791 -1189 1794 -1185
rect 1798 -1189 1808 -1185
rect 1791 -1191 1808 -1189
rect 1276 -1213 1282 -1211
rect 1276 -1217 1277 -1213
rect 1281 -1217 1282 -1213
rect 1276 -1219 1282 -1217
rect 1286 -1213 1303 -1211
rect 1286 -1217 1287 -1213
rect 1291 -1217 1303 -1213
rect 1286 -1219 1303 -1217
rect 1307 -1213 1324 -1211
rect 1307 -1217 1310 -1213
rect 1314 -1217 1324 -1213
rect 1307 -1219 1324 -1217
rect 946 -1232 963 -1230
rect 722 -1237 725 -1233
rect 729 -1237 739 -1233
rect 722 -1239 739 -1237
rect -107 -1277 -90 -1275
rect -578 -1279 -572 -1277
rect -578 -1283 -577 -1279
rect -573 -1283 -572 -1279
rect -578 -1285 -572 -1283
rect -568 -1279 -551 -1277
rect -568 -1283 -567 -1279
rect -563 -1283 -551 -1279
rect -568 -1285 -551 -1283
rect -547 -1279 -530 -1277
rect -547 -1283 -544 -1279
rect -540 -1283 -530 -1279
rect -547 -1285 -530 -1283
rect -512 -1279 -506 -1277
rect -512 -1283 -511 -1279
rect -507 -1283 -506 -1279
rect -512 -1285 -506 -1283
rect -502 -1279 -496 -1277
rect -502 -1283 -501 -1279
rect -497 -1283 -496 -1279
rect -502 -1285 -496 -1283
rect 605 -1274 611 -1272
rect 605 -1278 606 -1274
rect 610 -1278 611 -1274
rect 605 -1280 611 -1278
rect 615 -1274 632 -1272
rect 615 -1278 616 -1274
rect 620 -1278 632 -1274
rect 615 -1280 632 -1278
rect 636 -1274 653 -1272
rect 636 -1278 639 -1274
rect 643 -1278 653 -1274
rect 1674 -1226 1680 -1224
rect 1674 -1230 1675 -1226
rect 1679 -1230 1680 -1226
rect 1450 -1233 1456 -1231
rect 1450 -1237 1451 -1233
rect 1455 -1237 1456 -1233
rect 1450 -1239 1456 -1237
rect 1460 -1233 1477 -1231
rect 1460 -1237 1461 -1233
rect 1465 -1237 1477 -1233
rect 1460 -1239 1477 -1237
rect 1481 -1233 1498 -1231
rect 1674 -1232 1680 -1230
rect 1684 -1226 1701 -1224
rect 1684 -1230 1685 -1226
rect 1689 -1230 1701 -1226
rect 1684 -1232 1701 -1230
rect 1705 -1226 1722 -1224
rect 1705 -1230 1708 -1226
rect 1712 -1230 1722 -1226
rect 2496 -1185 2502 -1183
rect 2496 -1189 2497 -1185
rect 2501 -1189 2502 -1185
rect 2496 -1191 2502 -1189
rect 2506 -1185 2523 -1183
rect 2506 -1189 2507 -1185
rect 2511 -1189 2523 -1185
rect 2506 -1191 2523 -1189
rect 2527 -1185 2544 -1183
rect 2527 -1189 2530 -1185
rect 2534 -1189 2544 -1185
rect 2527 -1191 2544 -1189
rect 2012 -1213 2018 -1211
rect 2012 -1217 2013 -1213
rect 2017 -1217 2018 -1213
rect 2012 -1219 2018 -1217
rect 2022 -1213 2039 -1211
rect 2022 -1217 2023 -1213
rect 2027 -1217 2039 -1213
rect 2022 -1219 2039 -1217
rect 2043 -1213 2060 -1211
rect 2043 -1217 2046 -1213
rect 2050 -1217 2060 -1213
rect 2043 -1219 2060 -1217
rect 1705 -1232 1722 -1230
rect 1481 -1237 1484 -1233
rect 1488 -1237 1498 -1233
rect 1481 -1239 1498 -1237
rect 636 -1280 653 -1278
rect 1364 -1274 1370 -1272
rect 1364 -1278 1365 -1274
rect 1369 -1278 1370 -1274
rect 1364 -1280 1370 -1278
rect 1374 -1274 1391 -1272
rect 1374 -1278 1375 -1274
rect 1379 -1278 1391 -1274
rect 1374 -1280 1391 -1278
rect 1395 -1274 1412 -1272
rect 1395 -1278 1398 -1274
rect 1402 -1278 1412 -1274
rect 2410 -1226 2416 -1224
rect 2410 -1230 2411 -1226
rect 2415 -1230 2416 -1226
rect 2186 -1233 2192 -1231
rect 2186 -1237 2187 -1233
rect 2191 -1237 2192 -1233
rect 2186 -1239 2192 -1237
rect 2196 -1233 2213 -1231
rect 2196 -1237 2197 -1233
rect 2201 -1237 2213 -1233
rect 2196 -1239 2213 -1237
rect 2217 -1233 2234 -1231
rect 2410 -1232 2416 -1230
rect 2420 -1226 2437 -1224
rect 2420 -1230 2421 -1226
rect 2425 -1230 2437 -1226
rect 2420 -1232 2437 -1230
rect 2441 -1226 2458 -1224
rect 2441 -1230 2444 -1226
rect 2448 -1230 2458 -1226
rect 2441 -1232 2458 -1230
rect 2217 -1237 2220 -1233
rect 2224 -1237 2234 -1233
rect 2217 -1239 2234 -1237
rect 1395 -1280 1412 -1278
rect 2100 -1274 2106 -1272
rect 2100 -1278 2101 -1274
rect 2105 -1278 2106 -1274
rect 2100 -1280 2106 -1278
rect 2110 -1274 2127 -1272
rect 2110 -1278 2111 -1274
rect 2115 -1278 2127 -1274
rect 2110 -1280 2127 -1278
rect 2131 -1274 2148 -1272
rect 2131 -1278 2134 -1274
rect 2138 -1278 2148 -1274
rect 2131 -1280 2148 -1278
rect 144 -1329 150 -1327
rect 144 -1333 145 -1329
rect 149 -1333 150 -1329
rect 144 -1335 150 -1333
rect 154 -1329 171 -1327
rect 154 -1333 155 -1329
rect 159 -1333 171 -1329
rect 154 -1335 171 -1333
rect 175 -1329 192 -1327
rect 175 -1333 178 -1329
rect 182 -1333 192 -1329
rect 175 -1335 192 -1333
rect 210 -1329 216 -1327
rect 210 -1333 211 -1329
rect 215 -1333 216 -1329
rect 210 -1335 216 -1333
rect 220 -1329 226 -1327
rect 220 -1333 221 -1329
rect 225 -1333 226 -1329
rect 220 -1335 226 -1333
rect 303 -1329 309 -1327
rect 303 -1333 304 -1329
rect 308 -1333 309 -1329
rect 303 -1335 309 -1333
rect 313 -1335 330 -1327
rect 334 -1329 351 -1327
rect 334 -1333 339 -1329
rect 343 -1333 351 -1329
rect 334 -1335 351 -1333
rect 371 -1329 377 -1327
rect 371 -1333 372 -1329
rect 376 -1333 377 -1329
rect 371 -1335 377 -1333
rect 381 -1329 387 -1327
rect 381 -1333 382 -1329
rect 386 -1333 387 -1329
rect 887 -1332 893 -1330
rect 381 -1335 387 -1333
rect -581 -1371 -575 -1369
rect -581 -1375 -580 -1371
rect -576 -1375 -575 -1371
rect -581 -1377 -575 -1375
rect -571 -1371 -554 -1369
rect -571 -1375 -570 -1371
rect -566 -1375 -554 -1371
rect -571 -1377 -554 -1375
rect -550 -1371 -533 -1369
rect -550 -1375 -547 -1371
rect -543 -1375 -533 -1371
rect -550 -1377 -533 -1375
rect -515 -1371 -509 -1369
rect -515 -1375 -514 -1371
rect -510 -1375 -509 -1371
rect -515 -1377 -509 -1375
rect -505 -1371 -499 -1369
rect -505 -1375 -504 -1371
rect -500 -1375 -499 -1371
rect -505 -1377 -499 -1375
rect -167 -1380 -161 -1378
rect -167 -1384 -166 -1380
rect -162 -1384 -161 -1380
rect -167 -1386 -161 -1384
rect -157 -1380 -140 -1378
rect -157 -1384 -156 -1380
rect -152 -1384 -140 -1380
rect -157 -1386 -140 -1384
rect -136 -1380 -119 -1378
rect -136 -1384 -133 -1380
rect -129 -1384 -119 -1380
rect -136 -1386 -119 -1384
rect -101 -1380 -95 -1378
rect -101 -1384 -100 -1380
rect -96 -1384 -95 -1380
rect -101 -1386 -95 -1384
rect -91 -1380 -85 -1378
rect 887 -1336 888 -1332
rect 892 -1336 893 -1332
rect 887 -1338 893 -1336
rect 897 -1332 914 -1330
rect 897 -1336 898 -1332
rect 902 -1336 914 -1332
rect 897 -1338 914 -1336
rect 918 -1332 935 -1330
rect 918 -1336 921 -1332
rect 925 -1336 935 -1332
rect 918 -1338 935 -1336
rect 953 -1332 959 -1330
rect 953 -1336 954 -1332
rect 958 -1336 959 -1332
rect 953 -1338 959 -1336
rect 963 -1332 969 -1330
rect 963 -1336 964 -1332
rect 968 -1336 969 -1332
rect 963 -1338 969 -1336
rect 1046 -1332 1052 -1330
rect 1046 -1336 1047 -1332
rect 1051 -1336 1052 -1332
rect 1046 -1338 1052 -1336
rect 1056 -1338 1073 -1330
rect 1077 -1332 1094 -1330
rect 1077 -1336 1082 -1332
rect 1086 -1336 1094 -1332
rect 1077 -1338 1094 -1336
rect 1114 -1332 1120 -1330
rect 1114 -1336 1115 -1332
rect 1119 -1336 1120 -1332
rect 1114 -1338 1120 -1336
rect 1124 -1332 1130 -1330
rect 1124 -1336 1125 -1332
rect 1129 -1336 1130 -1332
rect 1646 -1332 1652 -1330
rect 1124 -1338 1130 -1336
rect 1646 -1336 1647 -1332
rect 1651 -1336 1652 -1332
rect 1646 -1338 1652 -1336
rect 1656 -1332 1673 -1330
rect 1656 -1336 1657 -1332
rect 1661 -1336 1673 -1332
rect 1656 -1338 1673 -1336
rect 1677 -1332 1694 -1330
rect 1677 -1336 1680 -1332
rect 1684 -1336 1694 -1332
rect 1677 -1338 1694 -1336
rect 1712 -1332 1718 -1330
rect 1712 -1336 1713 -1332
rect 1717 -1336 1718 -1332
rect 1712 -1338 1718 -1336
rect 1722 -1332 1728 -1330
rect 1722 -1336 1723 -1332
rect 1727 -1336 1728 -1332
rect 1722 -1338 1728 -1336
rect 1805 -1332 1811 -1330
rect 1805 -1336 1806 -1332
rect 1810 -1336 1811 -1332
rect 1805 -1338 1811 -1336
rect 1815 -1338 1832 -1330
rect 1836 -1332 1853 -1330
rect 1836 -1336 1841 -1332
rect 1845 -1336 1853 -1332
rect 1836 -1338 1853 -1336
rect 1873 -1332 1879 -1330
rect 1873 -1336 1874 -1332
rect 1878 -1336 1879 -1332
rect 1873 -1338 1879 -1336
rect 1883 -1332 1889 -1330
rect 1883 -1336 1884 -1332
rect 1888 -1336 1889 -1332
rect 2382 -1332 2388 -1330
rect 1883 -1338 1889 -1336
rect 2382 -1336 2383 -1332
rect 2387 -1336 2388 -1332
rect 2382 -1338 2388 -1336
rect 2392 -1332 2409 -1330
rect 2392 -1336 2393 -1332
rect 2397 -1336 2409 -1332
rect 2392 -1338 2409 -1336
rect 2413 -1332 2430 -1330
rect 2413 -1336 2416 -1332
rect 2420 -1336 2430 -1332
rect 2413 -1338 2430 -1336
rect 2448 -1332 2454 -1330
rect 2448 -1336 2449 -1332
rect 2453 -1336 2454 -1332
rect 2448 -1338 2454 -1336
rect 2458 -1332 2464 -1330
rect 2458 -1336 2459 -1332
rect 2463 -1336 2464 -1332
rect 2458 -1338 2464 -1336
rect 2541 -1332 2547 -1330
rect 2541 -1336 2542 -1332
rect 2546 -1336 2547 -1332
rect 2541 -1338 2547 -1336
rect 2551 -1338 2568 -1330
rect 2572 -1332 2589 -1330
rect 2572 -1336 2577 -1332
rect 2581 -1336 2589 -1332
rect 2572 -1338 2589 -1336
rect 2609 -1332 2615 -1330
rect 2609 -1336 2610 -1332
rect 2614 -1336 2615 -1332
rect 2609 -1338 2615 -1336
rect 2619 -1332 2625 -1330
rect 2619 -1336 2620 -1332
rect 2624 -1336 2625 -1332
rect 2619 -1338 2625 -1336
rect -91 -1384 -90 -1380
rect -86 -1384 -85 -1380
rect 576 -1383 582 -1381
rect -91 -1386 -85 -1384
rect 576 -1387 577 -1383
rect 581 -1387 582 -1383
rect 576 -1389 582 -1387
rect 586 -1383 603 -1381
rect 586 -1387 587 -1383
rect 591 -1387 603 -1383
rect 586 -1389 603 -1387
rect 607 -1383 624 -1381
rect 607 -1387 610 -1383
rect 614 -1387 624 -1383
rect 607 -1389 624 -1387
rect 642 -1383 648 -1381
rect 642 -1387 643 -1383
rect 647 -1387 648 -1383
rect 642 -1389 648 -1387
rect 652 -1383 658 -1381
rect 652 -1387 653 -1383
rect 657 -1387 658 -1383
rect 1335 -1383 1341 -1381
rect 652 -1389 658 -1387
rect 1335 -1387 1336 -1383
rect 1340 -1387 1341 -1383
rect 1335 -1389 1341 -1387
rect 1345 -1383 1362 -1381
rect 1345 -1387 1346 -1383
rect 1350 -1387 1362 -1383
rect 1345 -1389 1362 -1387
rect 1366 -1383 1383 -1381
rect 1366 -1387 1369 -1383
rect 1373 -1387 1383 -1383
rect 1366 -1389 1383 -1387
rect 1401 -1383 1407 -1381
rect 1401 -1387 1402 -1383
rect 1406 -1387 1407 -1383
rect 1401 -1389 1407 -1387
rect 1411 -1383 1417 -1381
rect 1411 -1387 1412 -1383
rect 1416 -1387 1417 -1383
rect 2071 -1383 2077 -1381
rect 1411 -1389 1417 -1387
rect 2071 -1387 2072 -1383
rect 2076 -1387 2077 -1383
rect 2071 -1389 2077 -1387
rect 2081 -1383 2098 -1381
rect 2081 -1387 2082 -1383
rect 2086 -1387 2098 -1383
rect 2081 -1389 2098 -1387
rect 2102 -1383 2119 -1381
rect 2102 -1387 2105 -1383
rect 2109 -1387 2119 -1383
rect 2102 -1389 2119 -1387
rect 2137 -1383 2143 -1381
rect 2137 -1387 2138 -1383
rect 2142 -1387 2143 -1383
rect 2137 -1389 2143 -1387
rect 2147 -1383 2153 -1381
rect 2147 -1387 2148 -1383
rect 2152 -1387 2153 -1383
rect 2147 -1389 2153 -1387
rect -581 -1463 -575 -1461
rect -581 -1467 -580 -1463
rect -576 -1467 -575 -1463
rect -581 -1469 -575 -1467
rect -571 -1463 -554 -1461
rect -571 -1467 -570 -1463
rect -566 -1467 -554 -1463
rect -571 -1469 -554 -1467
rect -550 -1463 -533 -1461
rect -550 -1467 -547 -1463
rect -543 -1467 -533 -1463
rect -550 -1469 -533 -1467
rect -515 -1463 -509 -1461
rect -515 -1467 -514 -1463
rect -510 -1467 -509 -1463
rect -515 -1469 -509 -1467
rect -505 -1463 -499 -1461
rect -505 -1467 -504 -1463
rect -500 -1467 -499 -1463
rect -505 -1469 -499 -1467
rect -581 -1555 -575 -1553
rect -581 -1559 -580 -1555
rect -576 -1559 -575 -1555
rect -581 -1561 -575 -1559
rect -571 -1555 -554 -1553
rect -571 -1559 -570 -1555
rect -566 -1559 -554 -1555
rect -571 -1561 -554 -1559
rect -550 -1555 -533 -1553
rect -550 -1559 -547 -1555
rect -543 -1559 -533 -1555
rect -550 -1561 -533 -1559
rect -515 -1555 -509 -1553
rect -515 -1559 -514 -1555
rect -510 -1559 -509 -1555
rect -515 -1561 -509 -1559
rect -505 -1555 -499 -1553
rect -505 -1559 -504 -1555
rect -500 -1559 -499 -1555
rect -505 -1561 -499 -1559
rect -580 -1675 -574 -1673
rect -580 -1679 -579 -1675
rect -575 -1679 -574 -1675
rect -580 -1681 -574 -1679
rect -570 -1675 -553 -1673
rect -570 -1679 -569 -1675
rect -565 -1679 -553 -1675
rect -570 -1681 -553 -1679
rect -549 -1675 -532 -1673
rect -549 -1679 -546 -1675
rect -542 -1679 -532 -1675
rect -549 -1681 -532 -1679
rect -514 -1675 -508 -1673
rect -514 -1679 -513 -1675
rect -509 -1679 -508 -1675
rect -514 -1681 -508 -1679
rect -504 -1675 -498 -1673
rect -504 -1679 -503 -1675
rect -499 -1679 -498 -1675
rect -504 -1681 -498 -1679
rect 13 -1731 19 -1729
rect 13 -1735 14 -1731
rect 18 -1735 19 -1731
rect 13 -1737 19 -1735
rect 23 -1731 40 -1729
rect 23 -1735 24 -1731
rect 28 -1735 40 -1731
rect 23 -1737 40 -1735
rect 44 -1731 61 -1729
rect 44 -1735 47 -1731
rect 51 -1735 61 -1731
rect 44 -1737 61 -1735
rect 502 -1731 508 -1729
rect 502 -1735 503 -1731
rect 507 -1735 508 -1731
rect 502 -1737 508 -1735
rect 512 -1731 529 -1729
rect 512 -1735 513 -1731
rect 517 -1735 529 -1731
rect 512 -1737 529 -1735
rect 533 -1731 550 -1729
rect 533 -1735 536 -1731
rect 540 -1735 550 -1731
rect 533 -1737 550 -1735
rect 886 -1731 892 -1729
rect 886 -1735 887 -1731
rect 891 -1735 892 -1731
rect 886 -1737 892 -1735
rect 896 -1731 913 -1729
rect 896 -1735 897 -1731
rect 901 -1735 913 -1731
rect 896 -1737 913 -1735
rect 917 -1731 934 -1729
rect 917 -1735 920 -1731
rect 924 -1735 934 -1731
rect 917 -1737 934 -1735
rect -583 -1767 -577 -1765
rect -583 -1771 -582 -1767
rect -578 -1771 -577 -1767
rect -583 -1773 -577 -1771
rect -573 -1767 -556 -1765
rect -573 -1771 -572 -1767
rect -568 -1771 -556 -1767
rect -573 -1773 -556 -1771
rect -552 -1767 -535 -1765
rect -552 -1771 -549 -1767
rect -545 -1771 -535 -1767
rect -552 -1773 -535 -1771
rect -517 -1767 -511 -1765
rect -517 -1771 -516 -1767
rect -512 -1771 -511 -1767
rect -517 -1773 -511 -1771
rect -507 -1767 -501 -1765
rect -507 -1771 -506 -1767
rect -502 -1771 -501 -1767
rect -507 -1773 -501 -1771
rect 1301 -1755 1307 -1753
rect 1301 -1759 1302 -1755
rect 1306 -1759 1307 -1755
rect 1301 -1761 1307 -1759
rect 1311 -1755 1328 -1753
rect 1311 -1759 1312 -1755
rect 1316 -1759 1328 -1755
rect 1311 -1761 1328 -1759
rect 1332 -1755 1349 -1753
rect 1332 -1759 1335 -1755
rect 1339 -1759 1349 -1755
rect 1332 -1761 1349 -1759
rect -60 -1779 -54 -1777
rect -60 -1783 -59 -1779
rect -55 -1783 -54 -1779
rect -60 -1785 -54 -1783
rect -50 -1779 -33 -1777
rect -50 -1783 -49 -1779
rect -45 -1783 -33 -1779
rect -50 -1785 -33 -1783
rect -29 -1779 -12 -1777
rect -29 -1783 -26 -1779
rect -22 -1783 -12 -1779
rect 429 -1779 435 -1777
rect -29 -1785 -12 -1783
rect 429 -1783 430 -1779
rect 434 -1783 435 -1779
rect 429 -1785 435 -1783
rect 439 -1779 456 -1777
rect 439 -1783 440 -1779
rect 444 -1783 456 -1779
rect 439 -1785 456 -1783
rect 460 -1779 477 -1777
rect 460 -1783 463 -1779
rect 467 -1783 477 -1779
rect 813 -1779 819 -1777
rect 460 -1785 477 -1783
rect 114 -1799 120 -1797
rect 114 -1803 115 -1799
rect 119 -1803 120 -1799
rect 114 -1805 120 -1803
rect 124 -1799 141 -1797
rect 124 -1803 125 -1799
rect 129 -1803 141 -1799
rect 124 -1805 141 -1803
rect 145 -1799 162 -1797
rect 145 -1803 148 -1799
rect 152 -1803 162 -1799
rect 145 -1805 162 -1803
rect 240 -1803 246 -1801
rect 28 -1840 34 -1838
rect 28 -1844 29 -1840
rect 33 -1844 34 -1840
rect 28 -1846 34 -1844
rect 38 -1840 55 -1838
rect 38 -1844 39 -1840
rect 43 -1844 55 -1840
rect 38 -1846 55 -1844
rect 59 -1840 76 -1838
rect 59 -1844 62 -1840
rect 66 -1844 76 -1840
rect 240 -1807 241 -1803
rect 245 -1807 246 -1803
rect 240 -1809 246 -1807
rect 250 -1803 256 -1801
rect 250 -1807 251 -1803
rect 255 -1807 256 -1803
rect 250 -1809 256 -1807
rect 813 -1783 814 -1779
rect 818 -1783 819 -1779
rect 813 -1785 819 -1783
rect 823 -1779 840 -1777
rect 823 -1783 824 -1779
rect 828 -1783 840 -1779
rect 823 -1785 840 -1783
rect 844 -1779 861 -1777
rect 844 -1783 847 -1779
rect 851 -1783 861 -1779
rect 844 -1785 861 -1783
rect 603 -1799 609 -1797
rect 603 -1803 604 -1799
rect 608 -1803 609 -1799
rect 603 -1805 609 -1803
rect 613 -1799 630 -1797
rect 613 -1803 614 -1799
rect 618 -1803 630 -1799
rect 613 -1805 630 -1803
rect 634 -1799 651 -1797
rect 634 -1803 637 -1799
rect 641 -1803 651 -1799
rect 634 -1805 651 -1803
rect 676 -1803 682 -1801
rect 517 -1840 523 -1838
rect 59 -1846 76 -1844
rect -583 -1859 -577 -1857
rect -583 -1863 -582 -1859
rect -578 -1863 -577 -1859
rect -583 -1865 -577 -1863
rect -573 -1859 -556 -1857
rect -573 -1863 -572 -1859
rect -568 -1863 -556 -1859
rect -573 -1865 -556 -1863
rect -552 -1859 -535 -1857
rect -552 -1863 -549 -1859
rect -545 -1863 -535 -1859
rect -552 -1865 -535 -1863
rect -517 -1859 -511 -1857
rect -517 -1863 -516 -1859
rect -512 -1863 -511 -1859
rect -517 -1865 -511 -1863
rect -507 -1859 -501 -1857
rect -507 -1863 -506 -1859
rect -502 -1863 -501 -1859
rect -507 -1865 -501 -1863
rect 517 -1844 518 -1840
rect 522 -1844 523 -1840
rect 517 -1846 523 -1844
rect 527 -1840 544 -1838
rect 527 -1844 528 -1840
rect 532 -1844 544 -1840
rect 527 -1846 544 -1844
rect 548 -1840 565 -1838
rect 548 -1844 551 -1840
rect 555 -1844 565 -1840
rect 676 -1807 677 -1803
rect 681 -1807 682 -1803
rect 676 -1809 682 -1807
rect 686 -1803 692 -1801
rect 686 -1807 687 -1803
rect 691 -1807 692 -1803
rect 686 -1809 692 -1807
rect 1021 -1799 1027 -1797
rect 1021 -1803 1022 -1799
rect 1026 -1803 1027 -1799
rect 1021 -1805 1027 -1803
rect 1031 -1799 1048 -1797
rect 1031 -1803 1032 -1799
rect 1036 -1803 1048 -1799
rect 1031 -1805 1048 -1803
rect 1052 -1799 1069 -1797
rect 1052 -1803 1055 -1799
rect 1059 -1803 1069 -1799
rect 1052 -1805 1069 -1803
rect 1094 -1803 1100 -1801
rect 901 -1840 907 -1838
rect 548 -1846 565 -1844
rect 901 -1844 902 -1840
rect 906 -1844 907 -1840
rect 901 -1846 907 -1844
rect 911 -1840 928 -1838
rect 911 -1844 912 -1840
rect 916 -1844 928 -1840
rect 911 -1846 928 -1844
rect 932 -1840 949 -1838
rect 932 -1844 935 -1840
rect 939 -1844 949 -1840
rect 1094 -1807 1095 -1803
rect 1099 -1807 1100 -1803
rect 1094 -1809 1100 -1807
rect 1104 -1803 1110 -1801
rect 1104 -1807 1105 -1803
rect 1109 -1807 1110 -1803
rect 1104 -1809 1110 -1807
rect 1228 -1803 1234 -1801
rect 1228 -1807 1229 -1803
rect 1233 -1807 1234 -1803
rect 1228 -1809 1234 -1807
rect 1238 -1803 1255 -1801
rect 1238 -1807 1239 -1803
rect 1243 -1807 1255 -1803
rect 1238 -1809 1255 -1807
rect 1259 -1803 1276 -1801
rect 1259 -1807 1262 -1803
rect 1266 -1807 1276 -1803
rect 1259 -1809 1276 -1807
rect 932 -1846 949 -1844
rect 1402 -1823 1408 -1821
rect 1402 -1827 1403 -1823
rect 1407 -1827 1408 -1823
rect 1402 -1829 1408 -1827
rect 1412 -1823 1429 -1821
rect 1412 -1827 1413 -1823
rect 1417 -1827 1429 -1823
rect 1412 -1829 1429 -1827
rect 1433 -1823 1450 -1821
rect 1433 -1827 1436 -1823
rect 1440 -1827 1450 -1823
rect 1433 -1829 1450 -1827
rect 1470 -1823 1476 -1821
rect 1470 -1827 1471 -1823
rect 1475 -1827 1476 -1823
rect 1470 -1829 1476 -1827
rect 1480 -1823 1486 -1821
rect 1480 -1827 1481 -1823
rect 1485 -1827 1486 -1823
rect 1480 -1829 1486 -1827
rect 1316 -1864 1322 -1862
rect 1316 -1868 1317 -1864
rect 1321 -1868 1322 -1864
rect 1316 -1870 1322 -1868
rect 1326 -1864 1343 -1862
rect 1326 -1868 1327 -1864
rect 1331 -1868 1343 -1864
rect 1326 -1870 1343 -1868
rect 1347 -1864 1364 -1862
rect 1347 -1868 1350 -1864
rect 1354 -1868 1364 -1864
rect 1347 -1870 1364 -1868
rect -583 -1951 -577 -1949
rect -583 -1955 -582 -1951
rect -578 -1955 -577 -1951
rect -583 -1957 -577 -1955
rect -573 -1951 -556 -1949
rect -573 -1955 -572 -1951
rect -568 -1955 -556 -1951
rect -573 -1957 -556 -1955
rect -552 -1951 -535 -1949
rect -552 -1955 -549 -1951
rect -545 -1955 -535 -1951
rect -552 -1957 -535 -1955
rect -517 -1951 -511 -1949
rect -517 -1955 -516 -1951
rect -512 -1955 -511 -1951
rect -517 -1957 -511 -1955
rect -507 -1951 -501 -1949
rect -507 -1955 -506 -1951
rect -502 -1955 -501 -1951
rect -507 -1957 -501 -1955
rect -578 -2042 -572 -2040
rect -578 -2046 -577 -2042
rect -573 -2046 -572 -2042
rect -578 -2048 -572 -2046
rect -568 -2042 -551 -2040
rect -568 -2046 -567 -2042
rect -563 -2046 -551 -2042
rect -568 -2048 -551 -2046
rect -547 -2042 -530 -2040
rect -547 -2046 -544 -2042
rect -540 -2046 -530 -2042
rect -547 -2048 -530 -2046
rect -512 -2042 -506 -2040
rect -512 -2046 -511 -2042
rect -507 -2046 -506 -2042
rect -512 -2048 -506 -2046
rect -502 -2042 -496 -2040
rect -502 -2046 -501 -2042
rect -497 -2046 -496 -2042
rect -502 -2048 -496 -2046
rect 333 -2089 339 -2087
rect 333 -2093 334 -2089
rect 338 -2093 339 -2089
rect 333 -2095 339 -2093
rect 343 -2089 372 -2087
rect 343 -2093 348 -2089
rect 352 -2093 372 -2089
rect 343 -2095 372 -2093
rect 376 -2089 396 -2087
rect 376 -2093 389 -2089
rect 393 -2093 396 -2089
rect 376 -2095 396 -2093
rect 400 -2089 418 -2087
rect 400 -2093 407 -2089
rect 411 -2093 418 -2089
rect 400 -2095 418 -2093
rect 441 -2089 447 -2087
rect 441 -2093 442 -2089
rect 446 -2093 447 -2089
rect 441 -2095 447 -2093
rect 451 -2089 457 -2087
rect 451 -2093 452 -2089
rect 456 -2093 457 -2089
rect 451 -2095 457 -2093
rect 749 -2089 755 -2087
rect 749 -2093 750 -2089
rect 754 -2093 755 -2089
rect 749 -2095 755 -2093
rect 759 -2089 788 -2087
rect 759 -2093 764 -2089
rect 768 -2093 788 -2089
rect 759 -2095 788 -2093
rect 792 -2089 812 -2087
rect 792 -2093 805 -2089
rect 809 -2093 812 -2089
rect 792 -2095 812 -2093
rect 816 -2089 834 -2087
rect 816 -2093 823 -2089
rect 827 -2093 834 -2089
rect 816 -2095 834 -2093
rect 857 -2089 863 -2087
rect 857 -2093 858 -2089
rect 862 -2093 863 -2089
rect 857 -2095 863 -2093
rect 867 -2089 873 -2087
rect 867 -2093 868 -2089
rect 872 -2093 873 -2089
rect 867 -2095 873 -2093
rect 1199 -2089 1205 -2087
rect 1199 -2093 1200 -2089
rect 1204 -2093 1205 -2089
rect 1199 -2095 1205 -2093
rect 1209 -2089 1238 -2087
rect 1209 -2093 1214 -2089
rect 1218 -2093 1238 -2089
rect 1209 -2095 1238 -2093
rect 1242 -2089 1262 -2087
rect 1242 -2093 1255 -2089
rect 1259 -2093 1262 -2089
rect 1242 -2095 1262 -2093
rect 1266 -2089 1284 -2087
rect 1266 -2093 1273 -2089
rect 1277 -2093 1284 -2089
rect 1266 -2095 1284 -2093
rect 1307 -2089 1313 -2087
rect 1307 -2093 1308 -2089
rect 1312 -2093 1313 -2089
rect 1307 -2095 1313 -2093
rect 1317 -2089 1323 -2087
rect 1317 -2093 1318 -2089
rect 1322 -2093 1323 -2089
rect 1317 -2095 1323 -2093
rect -581 -2134 -575 -2132
rect -581 -2138 -580 -2134
rect -576 -2138 -575 -2134
rect -581 -2140 -575 -2138
rect -571 -2134 -554 -2132
rect -571 -2138 -570 -2134
rect -566 -2138 -554 -2134
rect -571 -2140 -554 -2138
rect -550 -2134 -533 -2132
rect -550 -2138 -547 -2134
rect -543 -2138 -533 -2134
rect -550 -2140 -533 -2138
rect -515 -2134 -509 -2132
rect -515 -2138 -514 -2134
rect -510 -2138 -509 -2134
rect -515 -2140 -509 -2138
rect -505 -2134 -499 -2132
rect -505 -2138 -504 -2134
rect -500 -2138 -499 -2134
rect -505 -2140 -499 -2138
rect 255 -2142 261 -2140
rect 255 -2146 256 -2142
rect 260 -2146 261 -2142
rect 255 -2148 261 -2146
rect 265 -2142 271 -2140
rect 265 -2146 266 -2142
rect 270 -2146 271 -2142
rect 265 -2148 271 -2146
rect -34 -2166 -28 -2164
rect -34 -2170 -33 -2166
rect -29 -2170 -28 -2166
rect -34 -2172 -28 -2170
rect -24 -2166 -18 -2164
rect -24 -2170 -23 -2166
rect -19 -2170 -18 -2166
rect -24 -2172 -18 -2170
rect 53 -2174 59 -2172
rect 53 -2178 54 -2174
rect 58 -2178 59 -2174
rect 53 -2180 59 -2178
rect 63 -2174 80 -2172
rect 63 -2178 64 -2174
rect 68 -2178 80 -2174
rect 63 -2180 80 -2178
rect 84 -2174 101 -2172
rect 84 -2178 87 -2174
rect 91 -2178 101 -2174
rect 84 -2180 101 -2178
rect 119 -2174 125 -2172
rect 119 -2178 120 -2174
rect 124 -2178 125 -2174
rect 119 -2180 125 -2178
rect 129 -2174 135 -2172
rect 129 -2178 130 -2174
rect 134 -2178 135 -2174
rect 129 -2180 135 -2178
rect 671 -2142 677 -2140
rect 671 -2146 672 -2142
rect 676 -2146 677 -2142
rect 671 -2148 677 -2146
rect 681 -2142 687 -2140
rect 681 -2146 682 -2142
rect 686 -2146 687 -2142
rect 681 -2148 687 -2146
rect 1115 -2142 1121 -2140
rect 1115 -2146 1116 -2142
rect 1120 -2146 1121 -2142
rect 1115 -2148 1121 -2146
rect 1125 -2142 1131 -2140
rect 1125 -2146 1126 -2142
rect 1130 -2146 1131 -2142
rect 1125 -2148 1131 -2146
rect -581 -2226 -575 -2224
rect -581 -2230 -580 -2226
rect -576 -2230 -575 -2226
rect -581 -2232 -575 -2230
rect -571 -2226 -554 -2224
rect -571 -2230 -570 -2226
rect -566 -2230 -554 -2226
rect -571 -2232 -554 -2230
rect -550 -2226 -533 -2224
rect -550 -2230 -547 -2226
rect -543 -2230 -533 -2226
rect -550 -2232 -533 -2230
rect -515 -2226 -509 -2224
rect -515 -2230 -514 -2226
rect -510 -2230 -509 -2226
rect -515 -2232 -509 -2230
rect -505 -2226 -499 -2224
rect -505 -2230 -504 -2226
rect -500 -2230 -499 -2226
rect -505 -2232 -499 -2230
rect 351 -2226 357 -2224
rect 351 -2230 352 -2226
rect 356 -2230 357 -2226
rect 351 -2232 357 -2230
rect 361 -2226 390 -2224
rect 361 -2230 366 -2226
rect 370 -2230 390 -2226
rect 361 -2232 390 -2230
rect 394 -2226 414 -2224
rect 394 -2230 407 -2226
rect 411 -2230 414 -2226
rect 394 -2232 414 -2230
rect 418 -2226 436 -2224
rect 418 -2230 425 -2226
rect 429 -2230 436 -2226
rect 418 -2232 436 -2230
rect 459 -2226 465 -2224
rect 459 -2230 460 -2226
rect 464 -2230 465 -2226
rect 459 -2232 465 -2230
rect 469 -2226 475 -2224
rect 469 -2230 470 -2226
rect 474 -2230 475 -2226
rect 1217 -2226 1223 -2224
rect 469 -2232 475 -2230
rect 255 -2234 261 -2232
rect 255 -2238 256 -2234
rect 260 -2238 261 -2234
rect 255 -2240 261 -2238
rect 265 -2234 271 -2232
rect 265 -2238 266 -2234
rect 270 -2238 271 -2234
rect 265 -2240 271 -2238
rect -36 -2259 -30 -2257
rect -36 -2263 -35 -2259
rect -31 -2263 -30 -2259
rect -36 -2265 -30 -2263
rect -26 -2259 -20 -2257
rect -26 -2263 -25 -2259
rect -21 -2263 -20 -2259
rect -26 -2265 -20 -2263
rect 54 -2290 60 -2288
rect 54 -2294 55 -2290
rect 59 -2294 60 -2290
rect 54 -2296 60 -2294
rect 64 -2290 81 -2288
rect 64 -2294 65 -2290
rect 69 -2294 81 -2290
rect 64 -2296 81 -2294
rect 85 -2290 102 -2288
rect 85 -2294 88 -2290
rect 92 -2294 102 -2290
rect 85 -2296 102 -2294
rect 120 -2290 126 -2288
rect 120 -2294 121 -2290
rect 125 -2294 126 -2290
rect 120 -2296 126 -2294
rect 130 -2290 136 -2288
rect 130 -2294 131 -2290
rect 135 -2294 136 -2290
rect 130 -2296 136 -2294
rect -581 -2318 -575 -2316
rect -581 -2322 -580 -2318
rect -576 -2322 -575 -2318
rect -581 -2324 -575 -2322
rect -571 -2318 -554 -2316
rect -571 -2322 -570 -2318
rect -566 -2322 -554 -2318
rect -571 -2324 -554 -2322
rect -550 -2318 -533 -2316
rect -550 -2322 -547 -2318
rect -543 -2322 -533 -2318
rect -550 -2324 -533 -2322
rect -515 -2318 -509 -2316
rect -515 -2322 -514 -2318
rect -510 -2322 -509 -2318
rect -515 -2324 -509 -2322
rect -505 -2318 -499 -2316
rect -505 -2322 -504 -2318
rect -500 -2322 -499 -2318
rect -505 -2324 -499 -2322
rect 1217 -2230 1218 -2226
rect 1222 -2230 1223 -2226
rect 1217 -2232 1223 -2230
rect 1227 -2226 1256 -2224
rect 1227 -2230 1232 -2226
rect 1236 -2230 1256 -2226
rect 1227 -2232 1256 -2230
rect 1260 -2226 1280 -2224
rect 1260 -2230 1273 -2226
rect 1277 -2230 1280 -2226
rect 1260 -2232 1280 -2230
rect 1284 -2226 1302 -2224
rect 1284 -2230 1291 -2226
rect 1295 -2230 1302 -2226
rect 1284 -2232 1302 -2230
rect 1325 -2226 1331 -2224
rect 1325 -2230 1326 -2226
rect 1330 -2230 1331 -2226
rect 1325 -2232 1331 -2230
rect 1335 -2226 1341 -2224
rect 1335 -2230 1336 -2226
rect 1340 -2230 1341 -2226
rect 1335 -2232 1341 -2230
rect 1114 -2234 1120 -2232
rect 1114 -2238 1115 -2234
rect 1119 -2238 1120 -2234
rect 1114 -2240 1120 -2238
rect 1124 -2234 1130 -2232
rect 1124 -2238 1125 -2234
rect 1129 -2238 1130 -2234
rect 1124 -2240 1130 -2238
rect 767 -2254 773 -2252
rect 767 -2258 768 -2254
rect 772 -2258 773 -2254
rect 767 -2260 773 -2258
rect 777 -2254 806 -2252
rect 777 -2258 782 -2254
rect 786 -2258 806 -2254
rect 777 -2260 806 -2258
rect 810 -2254 830 -2252
rect 810 -2258 823 -2254
rect 827 -2258 830 -2254
rect 810 -2260 830 -2258
rect 834 -2254 852 -2252
rect 834 -2258 841 -2254
rect 845 -2258 852 -2254
rect 834 -2260 852 -2258
rect 875 -2254 881 -2252
rect 875 -2258 876 -2254
rect 880 -2258 881 -2254
rect 875 -2260 881 -2258
rect 885 -2254 891 -2252
rect 885 -2258 886 -2254
rect 890 -2258 891 -2254
rect 885 -2260 891 -2258
rect 664 -2262 670 -2260
rect 664 -2266 665 -2262
rect 669 -2266 670 -2262
rect 664 -2268 670 -2266
rect 674 -2262 680 -2260
rect 674 -2266 675 -2262
rect 679 -2266 680 -2262
rect 674 -2268 680 -2266
rect 547 -2311 553 -2309
rect 547 -2315 548 -2311
rect 552 -2315 553 -2311
rect 547 -2317 553 -2315
rect 557 -2311 574 -2309
rect 557 -2315 558 -2311
rect 562 -2315 574 -2311
rect 557 -2317 574 -2315
rect 578 -2311 595 -2309
rect 578 -2315 581 -2311
rect 585 -2315 595 -2311
rect 578 -2317 595 -2315
rect 613 -2311 619 -2309
rect 613 -2315 614 -2311
rect 618 -2315 619 -2311
rect 613 -2317 619 -2315
rect 623 -2311 629 -2309
rect 623 -2315 624 -2311
rect 628 -2315 629 -2311
rect 623 -2317 629 -2315
rect 956 -2272 962 -2270
rect 956 -2276 957 -2272
rect 961 -2276 962 -2272
rect 956 -2278 962 -2276
rect 966 -2272 983 -2270
rect 966 -2276 967 -2272
rect 971 -2276 983 -2272
rect 966 -2278 983 -2276
rect 987 -2272 1004 -2270
rect 987 -2276 990 -2272
rect 994 -2276 1004 -2272
rect 987 -2278 1004 -2276
rect 1022 -2272 1028 -2270
rect 1022 -2276 1023 -2272
rect 1027 -2276 1028 -2272
rect 1022 -2278 1028 -2276
rect 1032 -2272 1038 -2270
rect 1032 -2276 1033 -2272
rect 1037 -2276 1038 -2272
rect 1032 -2278 1038 -2276
rect 1437 -2267 1443 -2265
rect 1437 -2271 1438 -2267
rect 1442 -2271 1443 -2267
rect 1437 -2273 1443 -2271
rect 1447 -2267 1472 -2265
rect 1447 -2271 1448 -2267
rect 1452 -2271 1472 -2267
rect 1447 -2273 1472 -2271
rect 1476 -2267 1496 -2265
rect 1476 -2271 1489 -2267
rect 1493 -2271 1496 -2267
rect 1476 -2273 1496 -2271
rect 1500 -2267 1520 -2265
rect 1500 -2271 1509 -2267
rect 1513 -2271 1520 -2267
rect 1500 -2273 1520 -2271
rect 1524 -2267 1541 -2265
rect 1524 -2271 1530 -2267
rect 1534 -2271 1541 -2267
rect 1524 -2273 1541 -2271
rect 1561 -2267 1567 -2265
rect 1561 -2271 1562 -2267
rect 1566 -2271 1567 -2267
rect 1561 -2273 1567 -2271
rect 1571 -2267 1577 -2265
rect 1571 -2271 1572 -2267
rect 1576 -2271 1577 -2267
rect 1571 -2273 1577 -2271
rect 35 -2468 41 -2466
rect 35 -2472 36 -2468
rect 40 -2472 41 -2468
rect 35 -2474 41 -2472
rect 45 -2474 62 -2466
rect 66 -2474 83 -2466
rect 87 -2474 104 -2466
rect 108 -2468 146 -2466
rect 108 -2472 120 -2468
rect 124 -2472 146 -2468
rect 108 -2474 146 -2472
rect 166 -2468 172 -2466
rect 166 -2472 167 -2468
rect 171 -2472 172 -2468
rect 166 -2474 172 -2472
rect 176 -2468 182 -2466
rect 176 -2472 177 -2468
rect 181 -2472 182 -2468
rect 176 -2474 182 -2472
rect 305 -2468 311 -2466
rect 305 -2472 306 -2468
rect 310 -2472 311 -2468
rect 305 -2474 311 -2472
rect 315 -2474 332 -2466
rect 336 -2474 353 -2466
rect 357 -2474 374 -2466
rect 378 -2468 416 -2466
rect 378 -2472 390 -2468
rect 394 -2472 416 -2468
rect 378 -2474 416 -2472
rect 436 -2468 442 -2466
rect 436 -2472 437 -2468
rect 441 -2472 442 -2468
rect 436 -2474 442 -2472
rect 446 -2468 452 -2466
rect 446 -2472 447 -2468
rect 451 -2472 452 -2468
rect 446 -2474 452 -2472
rect -580 -2602 -574 -2600
rect -580 -2606 -579 -2602
rect -575 -2606 -574 -2602
rect -580 -2608 -574 -2606
rect -570 -2602 -553 -2600
rect -570 -2606 -569 -2602
rect -565 -2606 -553 -2602
rect -570 -2608 -553 -2606
rect -549 -2602 -532 -2600
rect -549 -2606 -546 -2602
rect -542 -2606 -532 -2602
rect -549 -2608 -532 -2606
rect -514 -2602 -508 -2600
rect -514 -2606 -513 -2602
rect -509 -2606 -508 -2602
rect -514 -2608 -508 -2606
rect -504 -2602 -498 -2600
rect -504 -2606 -503 -2602
rect -499 -2606 -498 -2602
rect -504 -2608 -498 -2606
rect -583 -2694 -577 -2692
rect -583 -2698 -582 -2694
rect -578 -2698 -577 -2694
rect -583 -2700 -577 -2698
rect -573 -2694 -556 -2692
rect -573 -2698 -572 -2694
rect -568 -2698 -556 -2694
rect -573 -2700 -556 -2698
rect -552 -2694 -535 -2692
rect -552 -2698 -549 -2694
rect -545 -2698 -535 -2694
rect -552 -2700 -535 -2698
rect -517 -2694 -511 -2692
rect -517 -2698 -516 -2694
rect -512 -2698 -511 -2694
rect -517 -2700 -511 -2698
rect -507 -2694 -501 -2692
rect -507 -2698 -506 -2694
rect -502 -2698 -501 -2694
rect -507 -2700 -501 -2698
rect -82 -2761 -76 -2759
rect -82 -2765 -81 -2761
rect -77 -2765 -76 -2761
rect -82 -2767 -76 -2765
rect -72 -2761 -55 -2759
rect -72 -2765 -71 -2761
rect -67 -2765 -55 -2761
rect -72 -2767 -55 -2765
rect -51 -2761 -34 -2759
rect -51 -2765 -48 -2761
rect -44 -2765 -34 -2761
rect -51 -2767 -34 -2765
rect -16 -2761 -10 -2759
rect -16 -2765 -15 -2761
rect -11 -2765 -10 -2761
rect -16 -2767 -10 -2765
rect -6 -2761 0 -2759
rect -6 -2765 -5 -2761
rect -1 -2765 0 -2761
rect -6 -2767 0 -2765
rect -583 -2786 -577 -2784
rect -583 -2790 -582 -2786
rect -578 -2790 -577 -2786
rect -583 -2792 -577 -2790
rect -573 -2786 -556 -2784
rect -573 -2790 -572 -2786
rect -568 -2790 -556 -2786
rect -573 -2792 -556 -2790
rect -552 -2786 -535 -2784
rect -552 -2790 -549 -2786
rect -545 -2790 -535 -2786
rect -552 -2792 -535 -2790
rect -517 -2786 -511 -2784
rect -517 -2790 -516 -2786
rect -512 -2790 -511 -2786
rect -517 -2792 -511 -2790
rect -507 -2786 -501 -2784
rect -507 -2790 -506 -2786
rect -502 -2790 -501 -2786
rect -507 -2792 -501 -2790
rect -82 -2854 -76 -2852
rect -82 -2858 -81 -2854
rect -77 -2858 -76 -2854
rect -82 -2860 -76 -2858
rect -72 -2854 -55 -2852
rect -72 -2858 -71 -2854
rect -67 -2858 -55 -2854
rect -72 -2860 -55 -2858
rect -51 -2854 -34 -2852
rect -51 -2858 -48 -2854
rect -44 -2858 -34 -2854
rect -51 -2860 -34 -2858
rect -16 -2854 -10 -2852
rect -16 -2858 -15 -2854
rect -11 -2858 -10 -2854
rect -16 -2860 -10 -2858
rect -6 -2854 0 -2852
rect -6 -2858 -5 -2854
rect -1 -2858 0 -2854
rect -6 -2860 0 -2858
rect -583 -2878 -577 -2876
rect -583 -2882 -582 -2878
rect -578 -2882 -577 -2878
rect -583 -2884 -577 -2882
rect -573 -2878 -556 -2876
rect -573 -2882 -572 -2878
rect -568 -2882 -556 -2878
rect -573 -2884 -556 -2882
rect -552 -2878 -535 -2876
rect -552 -2882 -549 -2878
rect -545 -2882 -535 -2878
rect -552 -2884 -535 -2882
rect -517 -2878 -511 -2876
rect -517 -2882 -516 -2878
rect -512 -2882 -511 -2878
rect -517 -2884 -511 -2882
rect -507 -2878 -501 -2876
rect -507 -2882 -506 -2878
rect -502 -2882 -501 -2878
rect -507 -2884 -501 -2882
rect -82 -2946 -76 -2944
rect -82 -2950 -81 -2946
rect -77 -2950 -76 -2946
rect -82 -2952 -76 -2950
rect -72 -2946 -55 -2944
rect -72 -2950 -71 -2946
rect -67 -2950 -55 -2946
rect -72 -2952 -55 -2950
rect -51 -2946 -34 -2944
rect -51 -2950 -48 -2946
rect -44 -2950 -34 -2946
rect -51 -2952 -34 -2950
rect -16 -2946 -10 -2944
rect -16 -2950 -15 -2946
rect -11 -2950 -10 -2946
rect -16 -2952 -10 -2950
rect -6 -2946 0 -2944
rect -6 -2950 -5 -2946
rect -1 -2950 0 -2946
rect -6 -2952 0 -2950
rect -578 -2969 -572 -2967
rect -578 -2973 -577 -2969
rect -573 -2973 -572 -2969
rect -578 -2975 -572 -2973
rect -568 -2969 -551 -2967
rect -568 -2973 -567 -2969
rect -563 -2973 -551 -2969
rect -568 -2975 -551 -2973
rect -547 -2969 -530 -2967
rect -547 -2973 -544 -2969
rect -540 -2973 -530 -2969
rect -547 -2975 -530 -2973
rect -512 -2969 -506 -2967
rect -512 -2973 -511 -2969
rect -507 -2973 -506 -2969
rect -512 -2975 -506 -2973
rect -502 -2969 -496 -2967
rect -502 -2973 -501 -2969
rect -497 -2973 -496 -2969
rect -502 -2975 -496 -2973
rect -82 -3039 -76 -3037
rect -82 -3043 -81 -3039
rect -77 -3043 -76 -3039
rect -82 -3045 -76 -3043
rect -72 -3039 -55 -3037
rect -72 -3043 -71 -3039
rect -67 -3043 -55 -3039
rect -72 -3045 -55 -3043
rect -51 -3039 -34 -3037
rect -51 -3043 -48 -3039
rect -44 -3043 -34 -3039
rect -51 -3045 -34 -3043
rect -16 -3039 -10 -3037
rect -16 -3043 -15 -3039
rect -11 -3043 -10 -3039
rect -16 -3045 -10 -3043
rect -6 -3039 0 -3037
rect -6 -3043 -5 -3039
rect -1 -3043 0 -3039
rect -6 -3045 0 -3043
rect -581 -3061 -575 -3059
rect -581 -3065 -580 -3061
rect -576 -3065 -575 -3061
rect -581 -3067 -575 -3065
rect -571 -3061 -554 -3059
rect -571 -3065 -570 -3061
rect -566 -3065 -554 -3061
rect -571 -3067 -554 -3065
rect -550 -3061 -533 -3059
rect -550 -3065 -547 -3061
rect -543 -3065 -533 -3061
rect -550 -3067 -533 -3065
rect -515 -3061 -509 -3059
rect -515 -3065 -514 -3061
rect -510 -3065 -509 -3061
rect -515 -3067 -509 -3065
rect -505 -3061 -499 -3059
rect -505 -3065 -504 -3061
rect -500 -3065 -499 -3061
rect -505 -3067 -499 -3065
rect -581 -3153 -575 -3151
rect -581 -3157 -580 -3153
rect -576 -3157 -575 -3153
rect -581 -3159 -575 -3157
rect -571 -3153 -554 -3151
rect -571 -3157 -570 -3153
rect -566 -3157 -554 -3153
rect -571 -3159 -554 -3157
rect -550 -3153 -533 -3151
rect -550 -3157 -547 -3153
rect -543 -3157 -533 -3153
rect -550 -3159 -533 -3157
rect -515 -3153 -509 -3151
rect -515 -3157 -514 -3153
rect -510 -3157 -509 -3153
rect -515 -3159 -509 -3157
rect -505 -3153 -499 -3151
rect -505 -3157 -504 -3153
rect -500 -3157 -499 -3153
rect -505 -3159 -499 -3157
rect -581 -3245 -575 -3243
rect -581 -3249 -580 -3245
rect -576 -3249 -575 -3245
rect -581 -3251 -575 -3249
rect -571 -3245 -554 -3243
rect -571 -3249 -570 -3245
rect -566 -3249 -554 -3245
rect -571 -3251 -554 -3249
rect -550 -3245 -533 -3243
rect -550 -3249 -547 -3245
rect -543 -3249 -533 -3245
rect -550 -3251 -533 -3249
rect -515 -3245 -509 -3243
rect -515 -3249 -514 -3245
rect -510 -3249 -509 -3245
rect -515 -3251 -509 -3249
rect -505 -3245 -499 -3243
rect -505 -3249 -504 -3245
rect -500 -3249 -499 -3245
rect -505 -3251 -499 -3249
<< ndcontact >>
rect -877 102 -873 106
rect -867 102 -863 106
rect -801 96 -797 100
rect -768 96 -764 100
rect -735 96 -731 100
rect -725 96 -721 100
rect -631 96 -627 100
rect -598 96 -594 100
rect -565 96 -561 100
rect -555 96 -551 100
rect -874 -7 -870 -3
rect -864 -7 -860 -3
rect -801 -13 -797 -9
rect -768 -13 -764 -9
rect -735 -13 -731 -9
rect -725 -13 -721 -9
rect -635 -13 -631 -9
rect -602 -13 -598 -9
rect -569 -13 -565 -9
rect -559 -13 -555 -9
rect -441 -14 -437 -10
rect -431 -14 -427 -10
rect -152 -67 -148 -63
rect -119 -67 -115 -63
rect 446 -67 450 -63
rect 479 -67 483 -63
rect -225 -115 -221 -111
rect -192 -115 -188 -111
rect 1325 -67 1329 -63
rect 1358 -67 1362 -63
rect 373 -115 377 -111
rect 406 -115 410 -111
rect -579 -168 -575 -164
rect -546 -168 -542 -164
rect -513 -168 -509 -164
rect -503 -168 -499 -164
rect -51 -135 -47 -131
rect -18 -135 -14 -131
rect 2093 -67 2097 -63
rect 2126 -67 2130 -63
rect 1252 -115 1256 -111
rect 1285 -115 1289 -111
rect 547 -135 551 -131
rect 580 -135 584 -131
rect 2020 -115 2024 -111
rect 2053 -115 2057 -111
rect 1426 -135 1430 -131
rect 1459 -135 1463 -131
rect 2194 -135 2198 -131
rect 2227 -135 2231 -131
rect -137 -176 -133 -172
rect -104 -176 -100 -172
rect 461 -176 465 -172
rect 494 -176 498 -172
rect 1340 -176 1344 -172
rect 1373 -176 1377 -172
rect 2108 -176 2112 -172
rect 2141 -176 2145 -172
rect -582 -260 -578 -256
rect -549 -260 -545 -256
rect -516 -260 -512 -256
rect -506 -260 -502 -256
rect -582 -352 -578 -348
rect -549 -352 -545 -348
rect -516 -352 -512 -348
rect -506 -352 -502 -348
rect 129 -370 133 -366
rect 162 -370 166 -366
rect 872 -373 876 -369
rect 905 -373 909 -369
rect -181 -418 -177 -414
rect -148 -418 -144 -414
rect 56 -418 60 -414
rect 89 -418 93 -414
rect -582 -444 -578 -440
rect -549 -444 -545 -440
rect -516 -444 -512 -440
rect -506 -444 -502 -440
rect 1631 -373 1635 -369
rect 1664 -373 1668 -369
rect 562 -421 566 -417
rect 595 -421 599 -417
rect 799 -421 803 -417
rect 832 -421 836 -417
rect -254 -466 -250 -462
rect -221 -466 -217 -462
rect 230 -438 234 -434
rect 263 -438 267 -434
rect 2367 -373 2371 -369
rect 2400 -373 2404 -369
rect 1321 -421 1325 -417
rect 1354 -421 1358 -417
rect 1558 -421 1562 -417
rect 1591 -421 1595 -417
rect 489 -469 493 -465
rect 522 -469 526 -465
rect 144 -479 148 -475
rect -80 -486 -76 -482
rect 177 -479 181 -475
rect -47 -486 -43 -482
rect 973 -441 977 -437
rect 1006 -441 1010 -437
rect 2057 -421 2061 -417
rect 2090 -421 2094 -417
rect 2294 -421 2298 -417
rect 2327 -421 2331 -417
rect 1248 -469 1252 -465
rect 1281 -469 1285 -465
rect 887 -482 891 -478
rect -166 -527 -162 -523
rect -133 -527 -129 -523
rect 663 -489 667 -485
rect 920 -482 924 -478
rect 696 -489 700 -485
rect 1732 -441 1736 -437
rect 1765 -441 1769 -437
rect 1984 -469 1988 -465
rect 2017 -469 2021 -465
rect 1646 -482 1650 -478
rect 1422 -489 1426 -485
rect 1679 -482 1683 -478
rect 1455 -489 1459 -485
rect 2468 -441 2472 -437
rect 2501 -441 2505 -437
rect 2382 -482 2386 -478
rect 2158 -489 2162 -485
rect 2415 -482 2419 -478
rect 2191 -489 2195 -485
rect -577 -535 -573 -531
rect -544 -535 -540 -531
rect -511 -535 -507 -531
rect -501 -535 -497 -531
rect 577 -530 581 -526
rect 610 -530 614 -526
rect 1336 -530 1340 -526
rect 1369 -530 1373 -526
rect 2072 -530 2076 -526
rect 2105 -530 2109 -526
rect 116 -585 120 -581
rect 149 -585 153 -581
rect 182 -585 186 -581
rect 192 -585 196 -581
rect 275 -588 279 -584
rect 285 -588 289 -584
rect 308 -588 312 -584
rect 343 -588 347 -584
rect 353 -588 357 -584
rect 859 -588 863 -584
rect -580 -627 -576 -623
rect -547 -627 -543 -623
rect -514 -627 -510 -623
rect -504 -627 -500 -623
rect 892 -588 896 -584
rect 925 -588 929 -584
rect 935 -588 939 -584
rect 1018 -591 1022 -587
rect 1028 -591 1032 -587
rect 1051 -591 1055 -587
rect 1086 -591 1090 -587
rect 1096 -591 1100 -587
rect 1618 -588 1622 -584
rect 1651 -588 1655 -584
rect 1684 -588 1688 -584
rect 1694 -588 1698 -584
rect 1777 -591 1781 -587
rect 1787 -591 1791 -587
rect 1810 -591 1814 -587
rect 1845 -591 1849 -587
rect 1855 -591 1859 -587
rect 2354 -588 2358 -584
rect 2387 -588 2391 -584
rect 2420 -588 2424 -584
rect 2430 -588 2434 -584
rect 2513 -591 2517 -587
rect 2523 -591 2527 -587
rect 2546 -591 2550 -587
rect 2581 -591 2585 -587
rect 2591 -591 2595 -587
rect -195 -636 -191 -632
rect -162 -636 -158 -632
rect -129 -636 -125 -632
rect -119 -636 -115 -632
rect 548 -639 552 -635
rect 581 -639 585 -635
rect 614 -639 618 -635
rect 624 -639 628 -635
rect 1307 -639 1311 -635
rect 1340 -639 1344 -635
rect 1373 -639 1377 -635
rect 1383 -639 1387 -635
rect 2043 -639 2047 -635
rect 2076 -639 2080 -635
rect 2109 -639 2113 -635
rect 2119 -639 2123 -635
rect -580 -719 -576 -715
rect -547 -719 -543 -715
rect -514 -719 -510 -715
rect -504 -719 -500 -715
rect -580 -811 -576 -807
rect -547 -811 -543 -807
rect -514 -811 -510 -807
rect -504 -811 -500 -807
rect -123 -860 -119 -856
rect -90 -860 -86 -856
rect 475 -860 479 -856
rect 508 -860 512 -856
rect -196 -908 -192 -904
rect -163 -908 -159 -904
rect 1354 -860 1358 -856
rect 1387 -860 1391 -856
rect 402 -908 406 -904
rect 435 -908 439 -904
rect -579 -961 -575 -957
rect -546 -961 -542 -957
rect -513 -961 -509 -957
rect -503 -961 -499 -957
rect -22 -928 -18 -924
rect 11 -928 15 -924
rect 2122 -860 2126 -856
rect 2155 -860 2159 -856
rect 1281 -908 1285 -904
rect 1314 -908 1318 -904
rect 576 -928 580 -924
rect 609 -928 613 -924
rect 2049 -908 2053 -904
rect 2082 -908 2086 -904
rect 1455 -928 1459 -924
rect 1488 -928 1492 -924
rect 2223 -928 2227 -924
rect 2256 -928 2260 -924
rect -108 -969 -104 -965
rect -75 -969 -71 -965
rect 490 -969 494 -965
rect 523 -969 527 -965
rect 1369 -969 1373 -965
rect 1402 -969 1406 -965
rect 2137 -969 2141 -965
rect 2170 -969 2174 -965
rect -582 -1053 -578 -1049
rect -549 -1053 -545 -1049
rect -516 -1053 -512 -1049
rect -506 -1053 -502 -1049
rect -582 -1145 -578 -1141
rect -549 -1145 -545 -1141
rect -516 -1145 -512 -1141
rect -506 -1145 -502 -1141
rect 158 -1163 162 -1159
rect 191 -1163 195 -1159
rect 901 -1166 905 -1162
rect 934 -1166 938 -1162
rect -152 -1211 -148 -1207
rect -119 -1211 -115 -1207
rect 85 -1211 89 -1207
rect 118 -1211 122 -1207
rect -582 -1237 -578 -1233
rect -549 -1237 -545 -1233
rect -516 -1237 -512 -1233
rect -506 -1237 -502 -1233
rect 1660 -1166 1664 -1162
rect 1693 -1166 1697 -1162
rect 591 -1214 595 -1210
rect 624 -1214 628 -1210
rect 828 -1214 832 -1210
rect 861 -1214 865 -1210
rect -225 -1259 -221 -1255
rect -192 -1259 -188 -1255
rect 259 -1231 263 -1227
rect 292 -1231 296 -1227
rect 2396 -1166 2400 -1162
rect 2429 -1166 2433 -1162
rect 1350 -1214 1354 -1210
rect 1383 -1214 1387 -1210
rect 1587 -1214 1591 -1210
rect 1620 -1214 1624 -1210
rect 518 -1262 522 -1258
rect 551 -1262 555 -1258
rect 173 -1272 177 -1268
rect -51 -1279 -47 -1275
rect 206 -1272 210 -1268
rect -18 -1279 -14 -1275
rect 1002 -1234 1006 -1230
rect 1035 -1234 1039 -1230
rect 2086 -1214 2090 -1210
rect 2119 -1214 2123 -1210
rect 2323 -1214 2327 -1210
rect 2356 -1214 2360 -1210
rect 1277 -1262 1281 -1258
rect 1310 -1262 1314 -1258
rect 916 -1275 920 -1271
rect -137 -1320 -133 -1316
rect -104 -1320 -100 -1316
rect 692 -1282 696 -1278
rect 949 -1275 953 -1271
rect 725 -1282 729 -1278
rect 1761 -1234 1765 -1230
rect 1794 -1234 1798 -1230
rect 2013 -1262 2017 -1258
rect 2046 -1262 2050 -1258
rect 1675 -1275 1679 -1271
rect 1451 -1282 1455 -1278
rect 1708 -1275 1712 -1271
rect 1484 -1282 1488 -1278
rect 2497 -1234 2501 -1230
rect 2530 -1234 2534 -1230
rect 2411 -1275 2415 -1271
rect 2187 -1282 2191 -1278
rect 2444 -1275 2448 -1271
rect 2220 -1282 2224 -1278
rect -577 -1328 -573 -1324
rect -544 -1328 -540 -1324
rect -511 -1328 -507 -1324
rect -501 -1328 -497 -1324
rect 606 -1323 610 -1319
rect 639 -1323 643 -1319
rect 1365 -1323 1369 -1319
rect 1398 -1323 1402 -1319
rect 2101 -1323 2105 -1319
rect 2134 -1323 2138 -1319
rect 145 -1378 149 -1374
rect 178 -1378 182 -1374
rect 211 -1378 215 -1374
rect 221 -1378 225 -1374
rect 304 -1381 308 -1377
rect 314 -1381 318 -1377
rect 337 -1381 341 -1377
rect 372 -1381 376 -1377
rect 382 -1381 386 -1377
rect 888 -1381 892 -1377
rect -580 -1420 -576 -1416
rect -547 -1420 -543 -1416
rect -514 -1420 -510 -1416
rect -504 -1420 -500 -1416
rect 921 -1381 925 -1377
rect 954 -1381 958 -1377
rect 964 -1381 968 -1377
rect 1047 -1384 1051 -1380
rect 1057 -1384 1061 -1380
rect 1080 -1384 1084 -1380
rect 1115 -1384 1119 -1380
rect 1125 -1384 1129 -1380
rect 1647 -1381 1651 -1377
rect 1680 -1381 1684 -1377
rect 1713 -1381 1717 -1377
rect 1723 -1381 1727 -1377
rect 1806 -1384 1810 -1380
rect 1816 -1384 1820 -1380
rect 1839 -1384 1843 -1380
rect 1874 -1384 1878 -1380
rect 1884 -1384 1888 -1380
rect 2383 -1381 2387 -1377
rect 2416 -1381 2420 -1377
rect 2449 -1381 2453 -1377
rect 2459 -1381 2463 -1377
rect 2542 -1384 2546 -1380
rect 2552 -1384 2556 -1380
rect 2575 -1384 2579 -1380
rect 2610 -1384 2614 -1380
rect 2620 -1384 2624 -1380
rect -166 -1429 -162 -1425
rect -133 -1429 -129 -1425
rect -100 -1429 -96 -1425
rect -90 -1429 -86 -1425
rect 577 -1432 581 -1428
rect 610 -1432 614 -1428
rect 643 -1432 647 -1428
rect 653 -1432 657 -1428
rect 1336 -1432 1340 -1428
rect 1369 -1432 1373 -1428
rect 1402 -1432 1406 -1428
rect 1412 -1432 1416 -1428
rect 2072 -1432 2076 -1428
rect 2105 -1432 2109 -1428
rect 2138 -1432 2142 -1428
rect 2148 -1432 2152 -1428
rect -580 -1512 -576 -1508
rect -547 -1512 -543 -1508
rect -514 -1512 -510 -1508
rect -504 -1512 -500 -1508
rect -580 -1604 -576 -1600
rect -547 -1604 -543 -1600
rect -514 -1604 -510 -1600
rect -504 -1604 -500 -1600
rect -579 -1724 -575 -1720
rect -546 -1724 -542 -1720
rect -513 -1724 -509 -1720
rect -503 -1724 -499 -1720
rect 14 -1780 18 -1776
rect 47 -1780 51 -1776
rect -582 -1816 -578 -1812
rect -549 -1816 -545 -1812
rect -516 -1816 -512 -1812
rect -506 -1816 -502 -1812
rect 503 -1780 507 -1776
rect 536 -1780 540 -1776
rect -59 -1828 -55 -1824
rect -26 -1828 -22 -1824
rect 887 -1780 891 -1776
rect 920 -1780 924 -1776
rect 430 -1828 434 -1824
rect 463 -1828 467 -1824
rect 115 -1848 119 -1844
rect 148 -1848 152 -1844
rect 241 -1846 245 -1842
rect 251 -1846 255 -1842
rect 814 -1828 818 -1824
rect 847 -1828 851 -1824
rect 604 -1848 608 -1844
rect 637 -1848 641 -1844
rect 677 -1846 681 -1842
rect 687 -1846 691 -1842
rect 1302 -1804 1306 -1800
rect 1335 -1804 1339 -1800
rect 1022 -1848 1026 -1844
rect 1055 -1848 1059 -1844
rect 1095 -1846 1099 -1842
rect 1105 -1846 1109 -1842
rect 1229 -1852 1233 -1848
rect 1262 -1852 1266 -1848
rect 1471 -1866 1475 -1862
rect 29 -1889 33 -1885
rect 62 -1889 66 -1885
rect 518 -1889 522 -1885
rect 551 -1889 555 -1885
rect 902 -1889 906 -1885
rect 935 -1889 939 -1885
rect -582 -1908 -578 -1904
rect -549 -1908 -545 -1904
rect -516 -1908 -512 -1904
rect -506 -1908 -502 -1904
rect 1403 -1872 1407 -1868
rect 1481 -1866 1485 -1862
rect 1436 -1872 1440 -1868
rect 1317 -1913 1321 -1909
rect 1350 -1913 1354 -1909
rect -582 -2000 -578 -1996
rect -549 -2000 -545 -1996
rect -516 -2000 -512 -1996
rect -506 -2000 -502 -1996
rect -577 -2091 -573 -2087
rect -544 -2091 -540 -2087
rect -511 -2091 -507 -2087
rect -501 -2091 -497 -2087
rect -580 -2183 -576 -2179
rect -547 -2183 -543 -2179
rect -514 -2183 -510 -2179
rect -504 -2183 -500 -2179
rect -33 -2209 -29 -2205
rect -23 -2209 -19 -2205
rect 334 -2167 338 -2163
rect 407 -2167 411 -2163
rect 442 -2167 446 -2163
rect 452 -2167 456 -2163
rect 750 -2167 754 -2163
rect 823 -2167 827 -2163
rect 858 -2167 862 -2163
rect 868 -2167 872 -2163
rect 1200 -2167 1204 -2163
rect 1273 -2167 1277 -2163
rect 1308 -2167 1312 -2163
rect 1318 -2167 1322 -2163
rect 256 -2191 260 -2187
rect 266 -2191 270 -2187
rect 672 -2191 676 -2187
rect 682 -2191 686 -2187
rect 1116 -2191 1120 -2187
rect 1126 -2191 1130 -2187
rect 54 -2223 58 -2219
rect 87 -2223 91 -2219
rect 120 -2223 124 -2219
rect 130 -2223 134 -2219
rect -580 -2275 -576 -2271
rect -547 -2275 -543 -2271
rect -514 -2275 -510 -2271
rect -504 -2275 -500 -2271
rect 256 -2283 260 -2279
rect 266 -2283 270 -2279
rect -35 -2302 -31 -2298
rect -25 -2302 -21 -2298
rect 352 -2304 356 -2300
rect 425 -2304 429 -2300
rect 460 -2304 464 -2300
rect 470 -2304 474 -2300
rect 665 -2311 669 -2307
rect 675 -2311 679 -2307
rect 55 -2339 59 -2335
rect 88 -2339 92 -2335
rect 121 -2339 125 -2335
rect 131 -2339 135 -2335
rect 1115 -2283 1119 -2279
rect 1125 -2283 1129 -2279
rect 1218 -2304 1222 -2300
rect 1291 -2304 1295 -2300
rect 1326 -2304 1330 -2300
rect 1336 -2304 1340 -2300
rect 957 -2321 961 -2317
rect 990 -2321 994 -2317
rect 1023 -2321 1027 -2317
rect 1033 -2321 1037 -2317
rect 768 -2332 772 -2328
rect 841 -2332 845 -2328
rect 876 -2332 880 -2328
rect 886 -2332 890 -2328
rect 1438 -2333 1442 -2329
rect 1530 -2333 1534 -2329
rect 1562 -2333 1566 -2329
rect 1572 -2333 1576 -2329
rect 548 -2360 552 -2356
rect -580 -2367 -576 -2363
rect -547 -2367 -543 -2363
rect -514 -2367 -510 -2363
rect 581 -2360 585 -2356
rect 614 -2360 618 -2356
rect 624 -2360 628 -2356
rect -504 -2367 -500 -2363
rect 36 -2540 40 -2536
rect 46 -2540 50 -2536
rect 69 -2540 73 -2536
rect 93 -2540 97 -2536
rect 167 -2540 171 -2536
rect 177 -2540 181 -2536
rect 306 -2543 310 -2539
rect 316 -2543 320 -2539
rect 339 -2543 343 -2539
rect 363 -2543 367 -2539
rect 437 -2543 441 -2539
rect 447 -2543 451 -2539
rect -579 -2651 -575 -2647
rect -546 -2651 -542 -2647
rect -513 -2651 -509 -2647
rect -503 -2651 -499 -2647
rect -582 -2743 -578 -2739
rect -549 -2743 -545 -2739
rect -516 -2743 -512 -2739
rect -506 -2743 -502 -2739
rect -81 -2810 -77 -2806
rect -48 -2810 -44 -2806
rect -15 -2810 -11 -2806
rect -5 -2810 -1 -2806
rect -582 -2835 -578 -2831
rect -549 -2835 -545 -2831
rect -516 -2835 -512 -2831
rect -506 -2835 -502 -2831
rect -81 -2903 -77 -2899
rect -48 -2903 -44 -2899
rect -15 -2903 -11 -2899
rect -5 -2903 -1 -2899
rect -582 -2927 -578 -2923
rect -549 -2927 -545 -2923
rect -516 -2927 -512 -2923
rect -506 -2927 -502 -2923
rect -81 -2995 -77 -2991
rect -48 -2995 -44 -2991
rect -15 -2995 -11 -2991
rect -5 -2995 -1 -2991
rect -577 -3018 -573 -3014
rect -544 -3018 -540 -3014
rect -511 -3018 -507 -3014
rect -501 -3018 -497 -3014
rect -81 -3088 -77 -3084
rect -48 -3088 -44 -3084
rect -15 -3088 -11 -3084
rect -5 -3088 -1 -3084
rect -580 -3110 -576 -3106
rect -547 -3110 -543 -3106
rect -514 -3110 -510 -3106
rect -504 -3110 -500 -3106
rect -580 -3202 -576 -3198
rect -547 -3202 -543 -3198
rect -514 -3202 -510 -3198
rect -504 -3202 -500 -3198
rect -580 -3294 -576 -3290
rect -547 -3294 -543 -3290
rect -514 -3294 -510 -3290
rect -504 -3294 -500 -3290
<< pdcontact >>
rect -877 141 -873 145
rect -867 141 -863 145
rect -801 141 -797 145
rect -791 141 -787 145
rect -768 141 -764 145
rect -735 141 -731 145
rect -725 141 -721 145
rect -631 141 -627 145
rect -621 141 -617 145
rect -598 141 -594 145
rect -565 141 -561 145
rect -555 141 -551 145
rect -874 32 -870 36
rect -864 32 -860 36
rect -801 32 -797 36
rect -791 32 -787 36
rect -768 32 -764 36
rect -735 32 -731 36
rect -725 32 -721 36
rect -635 32 -631 36
rect -625 32 -621 36
rect -602 32 -598 36
rect -569 32 -565 36
rect -559 32 -555 36
rect -441 32 -437 36
rect -431 32 -427 36
rect -152 -22 -148 -18
rect -142 -22 -138 -18
rect -119 -22 -115 -18
rect 446 -22 450 -18
rect 456 -22 460 -18
rect 479 -22 483 -18
rect 1325 -22 1329 -18
rect 1335 -22 1339 -18
rect 1358 -22 1362 -18
rect 2093 -22 2097 -18
rect 2103 -22 2107 -18
rect 2126 -22 2130 -18
rect -225 -70 -221 -66
rect -215 -70 -211 -66
rect -192 -70 -188 -66
rect 373 -70 377 -66
rect 383 -70 387 -66
rect 406 -70 410 -66
rect -51 -90 -47 -86
rect -41 -90 -37 -86
rect -18 -90 -14 -86
rect -579 -123 -575 -119
rect -569 -123 -565 -119
rect -546 -123 -542 -119
rect -513 -123 -509 -119
rect -503 -123 -499 -119
rect -137 -131 -133 -127
rect -127 -131 -123 -127
rect -104 -131 -100 -127
rect 1252 -70 1256 -66
rect 1262 -70 1266 -66
rect 1285 -70 1289 -66
rect 547 -90 551 -86
rect 557 -90 561 -86
rect 580 -90 584 -86
rect 461 -131 465 -127
rect 471 -131 475 -127
rect 494 -131 498 -127
rect 2020 -70 2024 -66
rect 2030 -70 2034 -66
rect 2053 -70 2057 -66
rect 1426 -90 1430 -86
rect 1436 -90 1440 -86
rect 1459 -90 1463 -86
rect 1340 -131 1344 -127
rect 1350 -131 1354 -127
rect 1373 -131 1377 -127
rect 2194 -90 2198 -86
rect 2204 -90 2208 -86
rect 2227 -90 2231 -86
rect 2108 -131 2112 -127
rect 2118 -131 2122 -127
rect 2141 -131 2145 -127
rect -582 -215 -578 -211
rect -572 -215 -568 -211
rect -549 -215 -545 -211
rect -516 -215 -512 -211
rect -506 -215 -502 -211
rect -582 -307 -578 -303
rect -572 -307 -568 -303
rect -549 -307 -545 -303
rect -516 -307 -512 -303
rect -506 -307 -502 -303
rect 129 -325 133 -321
rect 139 -325 143 -321
rect 162 -325 166 -321
rect 872 -328 876 -324
rect 882 -328 886 -324
rect 905 -328 909 -324
rect 1631 -328 1635 -324
rect 1641 -328 1645 -324
rect 1664 -328 1668 -324
rect 2367 -328 2371 -324
rect 2377 -328 2381 -324
rect 2400 -328 2404 -324
rect -181 -373 -177 -369
rect -171 -373 -167 -369
rect -148 -373 -144 -369
rect 56 -373 60 -369
rect 66 -373 70 -369
rect 89 -373 93 -369
rect -582 -399 -578 -395
rect -572 -399 -568 -395
rect -549 -399 -545 -395
rect -516 -399 -512 -395
rect -506 -399 -502 -395
rect 562 -376 566 -372
rect 572 -376 576 -372
rect 595 -376 599 -372
rect 799 -376 803 -372
rect 809 -376 813 -372
rect 832 -376 836 -372
rect 230 -393 234 -389
rect 240 -393 244 -389
rect 263 -393 267 -389
rect -254 -421 -250 -417
rect -244 -421 -240 -417
rect -221 -421 -217 -417
rect 144 -434 148 -430
rect -80 -441 -76 -437
rect -70 -441 -66 -437
rect 154 -434 158 -430
rect 177 -434 181 -430
rect 1321 -376 1325 -372
rect 1331 -376 1335 -372
rect 1354 -376 1358 -372
rect 1558 -376 1562 -372
rect 1568 -376 1572 -372
rect 1591 -376 1595 -372
rect 973 -396 977 -392
rect 983 -396 987 -392
rect 1006 -396 1010 -392
rect 489 -424 493 -420
rect 499 -424 503 -420
rect 522 -424 526 -420
rect -47 -441 -43 -437
rect -166 -482 -162 -478
rect -156 -482 -152 -478
rect -133 -482 -129 -478
rect 887 -437 891 -433
rect 663 -444 667 -440
rect 673 -444 677 -440
rect 897 -437 901 -433
rect 920 -437 924 -433
rect 2057 -376 2061 -372
rect 2067 -376 2071 -372
rect 2090 -376 2094 -372
rect 2294 -376 2298 -372
rect 2304 -376 2308 -372
rect 2327 -376 2331 -372
rect 1732 -396 1736 -392
rect 1742 -396 1746 -392
rect 1765 -396 1769 -392
rect 1248 -424 1252 -420
rect 1258 -424 1262 -420
rect 1281 -424 1285 -420
rect 696 -444 700 -440
rect -577 -490 -573 -486
rect -567 -490 -563 -486
rect -544 -490 -540 -486
rect -511 -490 -507 -486
rect -501 -490 -497 -486
rect 577 -485 581 -481
rect 587 -485 591 -481
rect 610 -485 614 -481
rect 1646 -437 1650 -433
rect 1422 -444 1426 -440
rect 1432 -444 1436 -440
rect 1656 -437 1660 -433
rect 1679 -437 1683 -433
rect 2468 -396 2472 -392
rect 2478 -396 2482 -392
rect 2501 -396 2505 -392
rect 1984 -424 1988 -420
rect 1994 -424 1998 -420
rect 2017 -424 2021 -420
rect 1455 -444 1459 -440
rect 1336 -485 1340 -481
rect 1346 -485 1350 -481
rect 1369 -485 1373 -481
rect 2382 -437 2386 -433
rect 2158 -444 2162 -440
rect 2168 -444 2172 -440
rect 2392 -437 2396 -433
rect 2415 -437 2419 -433
rect 2191 -444 2195 -440
rect 2072 -485 2076 -481
rect 2082 -485 2086 -481
rect 2105 -485 2109 -481
rect 116 -540 120 -536
rect 126 -540 130 -536
rect 149 -540 153 -536
rect 182 -540 186 -536
rect 192 -540 196 -536
rect 275 -540 279 -536
rect 310 -540 314 -536
rect 343 -540 347 -536
rect 353 -540 357 -536
rect -580 -582 -576 -578
rect -570 -582 -566 -578
rect -547 -582 -543 -578
rect -514 -582 -510 -578
rect -504 -582 -500 -578
rect -195 -591 -191 -587
rect -185 -591 -181 -587
rect -162 -591 -158 -587
rect -129 -591 -125 -587
rect 859 -543 863 -539
rect 869 -543 873 -539
rect 892 -543 896 -539
rect 925 -543 929 -539
rect 935 -543 939 -539
rect 1018 -543 1022 -539
rect 1053 -543 1057 -539
rect 1086 -543 1090 -539
rect 1096 -543 1100 -539
rect 1618 -543 1622 -539
rect 1628 -543 1632 -539
rect 1651 -543 1655 -539
rect 1684 -543 1688 -539
rect 1694 -543 1698 -539
rect 1777 -543 1781 -539
rect 1812 -543 1816 -539
rect 1845 -543 1849 -539
rect 1855 -543 1859 -539
rect 2354 -543 2358 -539
rect 2364 -543 2368 -539
rect 2387 -543 2391 -539
rect 2420 -543 2424 -539
rect 2430 -543 2434 -539
rect 2513 -543 2517 -539
rect 2548 -543 2552 -539
rect 2581 -543 2585 -539
rect 2591 -543 2595 -539
rect -119 -591 -115 -587
rect 548 -594 552 -590
rect 558 -594 562 -590
rect 581 -594 585 -590
rect 614 -594 618 -590
rect 624 -594 628 -590
rect 1307 -594 1311 -590
rect 1317 -594 1321 -590
rect 1340 -594 1344 -590
rect 1373 -594 1377 -590
rect 1383 -594 1387 -590
rect 2043 -594 2047 -590
rect 2053 -594 2057 -590
rect 2076 -594 2080 -590
rect 2109 -594 2113 -590
rect 2119 -594 2123 -590
rect -580 -674 -576 -670
rect -570 -674 -566 -670
rect -547 -674 -543 -670
rect -514 -674 -510 -670
rect -504 -674 -500 -670
rect -580 -766 -576 -762
rect -570 -766 -566 -762
rect -547 -766 -543 -762
rect -514 -766 -510 -762
rect -504 -766 -500 -762
rect -123 -815 -119 -811
rect -113 -815 -109 -811
rect -90 -815 -86 -811
rect 475 -815 479 -811
rect 485 -815 489 -811
rect 508 -815 512 -811
rect 1354 -815 1358 -811
rect 1364 -815 1368 -811
rect 1387 -815 1391 -811
rect 2122 -815 2126 -811
rect 2132 -815 2136 -811
rect 2155 -815 2159 -811
rect -196 -863 -192 -859
rect -186 -863 -182 -859
rect -163 -863 -159 -859
rect 402 -863 406 -859
rect 412 -863 416 -859
rect 435 -863 439 -859
rect -22 -883 -18 -879
rect -12 -883 -8 -879
rect 11 -883 15 -879
rect -579 -916 -575 -912
rect -569 -916 -565 -912
rect -546 -916 -542 -912
rect -513 -916 -509 -912
rect -503 -916 -499 -912
rect -108 -924 -104 -920
rect -98 -924 -94 -920
rect -75 -924 -71 -920
rect 1281 -863 1285 -859
rect 1291 -863 1295 -859
rect 1314 -863 1318 -859
rect 576 -883 580 -879
rect 586 -883 590 -879
rect 609 -883 613 -879
rect 490 -924 494 -920
rect 500 -924 504 -920
rect 523 -924 527 -920
rect 2049 -863 2053 -859
rect 2059 -863 2063 -859
rect 2082 -863 2086 -859
rect 1455 -883 1459 -879
rect 1465 -883 1469 -879
rect 1488 -883 1492 -879
rect 1369 -924 1373 -920
rect 1379 -924 1383 -920
rect 1402 -924 1406 -920
rect 2223 -883 2227 -879
rect 2233 -883 2237 -879
rect 2256 -883 2260 -879
rect 2137 -924 2141 -920
rect 2147 -924 2151 -920
rect 2170 -924 2174 -920
rect -582 -1008 -578 -1004
rect -572 -1008 -568 -1004
rect -549 -1008 -545 -1004
rect -516 -1008 -512 -1004
rect -506 -1008 -502 -1004
rect -582 -1100 -578 -1096
rect -572 -1100 -568 -1096
rect -549 -1100 -545 -1096
rect -516 -1100 -512 -1096
rect -506 -1100 -502 -1096
rect 158 -1118 162 -1114
rect 168 -1118 172 -1114
rect 191 -1118 195 -1114
rect 901 -1121 905 -1117
rect 911 -1121 915 -1117
rect 934 -1121 938 -1117
rect 1660 -1121 1664 -1117
rect 1670 -1121 1674 -1117
rect 1693 -1121 1697 -1117
rect 2396 -1121 2400 -1117
rect 2406 -1121 2410 -1117
rect 2429 -1121 2433 -1117
rect -152 -1166 -148 -1162
rect -142 -1166 -138 -1162
rect -119 -1166 -115 -1162
rect 85 -1166 89 -1162
rect 95 -1166 99 -1162
rect 118 -1166 122 -1162
rect -582 -1192 -578 -1188
rect -572 -1192 -568 -1188
rect -549 -1192 -545 -1188
rect -516 -1192 -512 -1188
rect -506 -1192 -502 -1188
rect 591 -1169 595 -1165
rect 601 -1169 605 -1165
rect 624 -1169 628 -1165
rect 828 -1169 832 -1165
rect 838 -1169 842 -1165
rect 861 -1169 865 -1165
rect 259 -1186 263 -1182
rect 269 -1186 273 -1182
rect 292 -1186 296 -1182
rect -225 -1214 -221 -1210
rect -215 -1214 -211 -1210
rect -192 -1214 -188 -1210
rect 173 -1227 177 -1223
rect -51 -1234 -47 -1230
rect -41 -1234 -37 -1230
rect 183 -1227 187 -1223
rect 206 -1227 210 -1223
rect 1350 -1169 1354 -1165
rect 1360 -1169 1364 -1165
rect 1383 -1169 1387 -1165
rect 1587 -1169 1591 -1165
rect 1597 -1169 1601 -1165
rect 1620 -1169 1624 -1165
rect 1002 -1189 1006 -1185
rect 1012 -1189 1016 -1185
rect 1035 -1189 1039 -1185
rect 518 -1217 522 -1213
rect 528 -1217 532 -1213
rect 551 -1217 555 -1213
rect -18 -1234 -14 -1230
rect -137 -1275 -133 -1271
rect -127 -1275 -123 -1271
rect -104 -1275 -100 -1271
rect 916 -1230 920 -1226
rect 692 -1237 696 -1233
rect 702 -1237 706 -1233
rect 926 -1230 930 -1226
rect 949 -1230 953 -1226
rect 2086 -1169 2090 -1165
rect 2096 -1169 2100 -1165
rect 2119 -1169 2123 -1165
rect 2323 -1169 2327 -1165
rect 2333 -1169 2337 -1165
rect 2356 -1169 2360 -1165
rect 1761 -1189 1765 -1185
rect 1771 -1189 1775 -1185
rect 1794 -1189 1798 -1185
rect 1277 -1217 1281 -1213
rect 1287 -1217 1291 -1213
rect 1310 -1217 1314 -1213
rect 725 -1237 729 -1233
rect -577 -1283 -573 -1279
rect -567 -1283 -563 -1279
rect -544 -1283 -540 -1279
rect -511 -1283 -507 -1279
rect -501 -1283 -497 -1279
rect 606 -1278 610 -1274
rect 616 -1278 620 -1274
rect 639 -1278 643 -1274
rect 1675 -1230 1679 -1226
rect 1451 -1237 1455 -1233
rect 1461 -1237 1465 -1233
rect 1685 -1230 1689 -1226
rect 1708 -1230 1712 -1226
rect 2497 -1189 2501 -1185
rect 2507 -1189 2511 -1185
rect 2530 -1189 2534 -1185
rect 2013 -1217 2017 -1213
rect 2023 -1217 2027 -1213
rect 2046 -1217 2050 -1213
rect 1484 -1237 1488 -1233
rect 1365 -1278 1369 -1274
rect 1375 -1278 1379 -1274
rect 1398 -1278 1402 -1274
rect 2411 -1230 2415 -1226
rect 2187 -1237 2191 -1233
rect 2197 -1237 2201 -1233
rect 2421 -1230 2425 -1226
rect 2444 -1230 2448 -1226
rect 2220 -1237 2224 -1233
rect 2101 -1278 2105 -1274
rect 2111 -1278 2115 -1274
rect 2134 -1278 2138 -1274
rect 145 -1333 149 -1329
rect 155 -1333 159 -1329
rect 178 -1333 182 -1329
rect 211 -1333 215 -1329
rect 221 -1333 225 -1329
rect 304 -1333 308 -1329
rect 339 -1333 343 -1329
rect 372 -1333 376 -1329
rect 382 -1333 386 -1329
rect -580 -1375 -576 -1371
rect -570 -1375 -566 -1371
rect -547 -1375 -543 -1371
rect -514 -1375 -510 -1371
rect -504 -1375 -500 -1371
rect -166 -1384 -162 -1380
rect -156 -1384 -152 -1380
rect -133 -1384 -129 -1380
rect -100 -1384 -96 -1380
rect 888 -1336 892 -1332
rect 898 -1336 902 -1332
rect 921 -1336 925 -1332
rect 954 -1336 958 -1332
rect 964 -1336 968 -1332
rect 1047 -1336 1051 -1332
rect 1082 -1336 1086 -1332
rect 1115 -1336 1119 -1332
rect 1125 -1336 1129 -1332
rect 1647 -1336 1651 -1332
rect 1657 -1336 1661 -1332
rect 1680 -1336 1684 -1332
rect 1713 -1336 1717 -1332
rect 1723 -1336 1727 -1332
rect 1806 -1336 1810 -1332
rect 1841 -1336 1845 -1332
rect 1874 -1336 1878 -1332
rect 1884 -1336 1888 -1332
rect 2383 -1336 2387 -1332
rect 2393 -1336 2397 -1332
rect 2416 -1336 2420 -1332
rect 2449 -1336 2453 -1332
rect 2459 -1336 2463 -1332
rect 2542 -1336 2546 -1332
rect 2577 -1336 2581 -1332
rect 2610 -1336 2614 -1332
rect 2620 -1336 2624 -1332
rect -90 -1384 -86 -1380
rect 577 -1387 581 -1383
rect 587 -1387 591 -1383
rect 610 -1387 614 -1383
rect 643 -1387 647 -1383
rect 653 -1387 657 -1383
rect 1336 -1387 1340 -1383
rect 1346 -1387 1350 -1383
rect 1369 -1387 1373 -1383
rect 1402 -1387 1406 -1383
rect 1412 -1387 1416 -1383
rect 2072 -1387 2076 -1383
rect 2082 -1387 2086 -1383
rect 2105 -1387 2109 -1383
rect 2138 -1387 2142 -1383
rect 2148 -1387 2152 -1383
rect -580 -1467 -576 -1463
rect -570 -1467 -566 -1463
rect -547 -1467 -543 -1463
rect -514 -1467 -510 -1463
rect -504 -1467 -500 -1463
rect -580 -1559 -576 -1555
rect -570 -1559 -566 -1555
rect -547 -1559 -543 -1555
rect -514 -1559 -510 -1555
rect -504 -1559 -500 -1555
rect -579 -1679 -575 -1675
rect -569 -1679 -565 -1675
rect -546 -1679 -542 -1675
rect -513 -1679 -509 -1675
rect -503 -1679 -499 -1675
rect 14 -1735 18 -1731
rect 24 -1735 28 -1731
rect 47 -1735 51 -1731
rect 503 -1735 507 -1731
rect 513 -1735 517 -1731
rect 536 -1735 540 -1731
rect 887 -1735 891 -1731
rect 897 -1735 901 -1731
rect 920 -1735 924 -1731
rect -582 -1771 -578 -1767
rect -572 -1771 -568 -1767
rect -549 -1771 -545 -1767
rect -516 -1771 -512 -1767
rect -506 -1771 -502 -1767
rect 1302 -1759 1306 -1755
rect 1312 -1759 1316 -1755
rect 1335 -1759 1339 -1755
rect -59 -1783 -55 -1779
rect -49 -1783 -45 -1779
rect -26 -1783 -22 -1779
rect 430 -1783 434 -1779
rect 440 -1783 444 -1779
rect 463 -1783 467 -1779
rect 115 -1803 119 -1799
rect 125 -1803 129 -1799
rect 148 -1803 152 -1799
rect 29 -1844 33 -1840
rect 39 -1844 43 -1840
rect 62 -1844 66 -1840
rect 241 -1807 245 -1803
rect 251 -1807 255 -1803
rect 814 -1783 818 -1779
rect 824 -1783 828 -1779
rect 847 -1783 851 -1779
rect 604 -1803 608 -1799
rect 614 -1803 618 -1799
rect 637 -1803 641 -1799
rect -582 -1863 -578 -1859
rect -572 -1863 -568 -1859
rect -549 -1863 -545 -1859
rect -516 -1863 -512 -1859
rect -506 -1863 -502 -1859
rect 518 -1844 522 -1840
rect 528 -1844 532 -1840
rect 551 -1844 555 -1840
rect 677 -1807 681 -1803
rect 687 -1807 691 -1803
rect 1022 -1803 1026 -1799
rect 1032 -1803 1036 -1799
rect 1055 -1803 1059 -1799
rect 902 -1844 906 -1840
rect 912 -1844 916 -1840
rect 935 -1844 939 -1840
rect 1095 -1807 1099 -1803
rect 1105 -1807 1109 -1803
rect 1229 -1807 1233 -1803
rect 1239 -1807 1243 -1803
rect 1262 -1807 1266 -1803
rect 1403 -1827 1407 -1823
rect 1413 -1827 1417 -1823
rect 1436 -1827 1440 -1823
rect 1471 -1827 1475 -1823
rect 1481 -1827 1485 -1823
rect 1317 -1868 1321 -1864
rect 1327 -1868 1331 -1864
rect 1350 -1868 1354 -1864
rect -582 -1955 -578 -1951
rect -572 -1955 -568 -1951
rect -549 -1955 -545 -1951
rect -516 -1955 -512 -1951
rect -506 -1955 -502 -1951
rect -577 -2046 -573 -2042
rect -567 -2046 -563 -2042
rect -544 -2046 -540 -2042
rect -511 -2046 -507 -2042
rect -501 -2046 -497 -2042
rect 334 -2093 338 -2089
rect 348 -2093 352 -2089
rect 389 -2093 393 -2089
rect 407 -2093 411 -2089
rect 442 -2093 446 -2089
rect 452 -2093 456 -2089
rect 750 -2093 754 -2089
rect 764 -2093 768 -2089
rect 805 -2093 809 -2089
rect 823 -2093 827 -2089
rect 858 -2093 862 -2089
rect 868 -2093 872 -2089
rect 1200 -2093 1204 -2089
rect 1214 -2093 1218 -2089
rect 1255 -2093 1259 -2089
rect 1273 -2093 1277 -2089
rect 1308 -2093 1312 -2089
rect 1318 -2093 1322 -2089
rect -580 -2138 -576 -2134
rect -570 -2138 -566 -2134
rect -547 -2138 -543 -2134
rect -514 -2138 -510 -2134
rect -504 -2138 -500 -2134
rect 256 -2146 260 -2142
rect 266 -2146 270 -2142
rect -33 -2170 -29 -2166
rect -23 -2170 -19 -2166
rect 54 -2178 58 -2174
rect 64 -2178 68 -2174
rect 87 -2178 91 -2174
rect 120 -2178 124 -2174
rect 130 -2178 134 -2174
rect 672 -2146 676 -2142
rect 682 -2146 686 -2142
rect 1116 -2146 1120 -2142
rect 1126 -2146 1130 -2142
rect -580 -2230 -576 -2226
rect -570 -2230 -566 -2226
rect -547 -2230 -543 -2226
rect -514 -2230 -510 -2226
rect -504 -2230 -500 -2226
rect 352 -2230 356 -2226
rect 366 -2230 370 -2226
rect 407 -2230 411 -2226
rect 425 -2230 429 -2226
rect 460 -2230 464 -2226
rect 470 -2230 474 -2226
rect 256 -2238 260 -2234
rect 266 -2238 270 -2234
rect -35 -2263 -31 -2259
rect -25 -2263 -21 -2259
rect 55 -2294 59 -2290
rect 65 -2294 69 -2290
rect 88 -2294 92 -2290
rect 121 -2294 125 -2290
rect 131 -2294 135 -2290
rect -580 -2322 -576 -2318
rect -570 -2322 -566 -2318
rect -547 -2322 -543 -2318
rect -514 -2322 -510 -2318
rect -504 -2322 -500 -2318
rect 1218 -2230 1222 -2226
rect 1232 -2230 1236 -2226
rect 1273 -2230 1277 -2226
rect 1291 -2230 1295 -2226
rect 1326 -2230 1330 -2226
rect 1336 -2230 1340 -2226
rect 1115 -2238 1119 -2234
rect 1125 -2238 1129 -2234
rect 768 -2258 772 -2254
rect 782 -2258 786 -2254
rect 823 -2258 827 -2254
rect 841 -2258 845 -2254
rect 876 -2258 880 -2254
rect 886 -2258 890 -2254
rect 665 -2266 669 -2262
rect 675 -2266 679 -2262
rect 548 -2315 552 -2311
rect 558 -2315 562 -2311
rect 581 -2315 585 -2311
rect 614 -2315 618 -2311
rect 624 -2315 628 -2311
rect 957 -2276 961 -2272
rect 967 -2276 971 -2272
rect 990 -2276 994 -2272
rect 1023 -2276 1027 -2272
rect 1033 -2276 1037 -2272
rect 1438 -2271 1442 -2267
rect 1448 -2271 1452 -2267
rect 1489 -2271 1493 -2267
rect 1509 -2271 1513 -2267
rect 1530 -2271 1534 -2267
rect 1562 -2271 1566 -2267
rect 1572 -2271 1576 -2267
rect 36 -2472 40 -2468
rect 120 -2472 124 -2468
rect 167 -2472 171 -2468
rect 177 -2472 181 -2468
rect 306 -2472 310 -2468
rect 390 -2472 394 -2468
rect 437 -2472 441 -2468
rect 447 -2472 451 -2468
rect -579 -2606 -575 -2602
rect -569 -2606 -565 -2602
rect -546 -2606 -542 -2602
rect -513 -2606 -509 -2602
rect -503 -2606 -499 -2602
rect -582 -2698 -578 -2694
rect -572 -2698 -568 -2694
rect -549 -2698 -545 -2694
rect -516 -2698 -512 -2694
rect -506 -2698 -502 -2694
rect -81 -2765 -77 -2761
rect -71 -2765 -67 -2761
rect -48 -2765 -44 -2761
rect -15 -2765 -11 -2761
rect -5 -2765 -1 -2761
rect -582 -2790 -578 -2786
rect -572 -2790 -568 -2786
rect -549 -2790 -545 -2786
rect -516 -2790 -512 -2786
rect -506 -2790 -502 -2786
rect -81 -2858 -77 -2854
rect -71 -2858 -67 -2854
rect -48 -2858 -44 -2854
rect -15 -2858 -11 -2854
rect -5 -2858 -1 -2854
rect -582 -2882 -578 -2878
rect -572 -2882 -568 -2878
rect -549 -2882 -545 -2878
rect -516 -2882 -512 -2878
rect -506 -2882 -502 -2878
rect -81 -2950 -77 -2946
rect -71 -2950 -67 -2946
rect -48 -2950 -44 -2946
rect -15 -2950 -11 -2946
rect -5 -2950 -1 -2946
rect -577 -2973 -573 -2969
rect -567 -2973 -563 -2969
rect -544 -2973 -540 -2969
rect -511 -2973 -507 -2969
rect -501 -2973 -497 -2969
rect -81 -3043 -77 -3039
rect -71 -3043 -67 -3039
rect -48 -3043 -44 -3039
rect -15 -3043 -11 -3039
rect -5 -3043 -1 -3039
rect -580 -3065 -576 -3061
rect -570 -3065 -566 -3061
rect -547 -3065 -543 -3061
rect -514 -3065 -510 -3061
rect -504 -3065 -500 -3061
rect -580 -3157 -576 -3153
rect -570 -3157 -566 -3153
rect -547 -3157 -543 -3153
rect -514 -3157 -510 -3153
rect -504 -3157 -500 -3153
rect -580 -3249 -576 -3245
rect -570 -3249 -566 -3245
rect -547 -3249 -543 -3245
rect -514 -3249 -510 -3245
rect -504 -3249 -500 -3245
<< polysilicon >>
rect -872 147 -868 150
rect -796 147 -792 150
rect -775 147 -771 150
rect -730 147 -726 150
rect -626 147 -622 150
rect -605 147 -601 150
rect -560 147 -556 150
rect -872 108 -868 139
rect -796 102 -792 139
rect -775 102 -771 139
rect -730 102 -726 139
rect -626 102 -622 139
rect -605 102 -601 139
rect -560 102 -556 139
rect -872 97 -868 100
rect -796 91 -792 94
rect -775 91 -771 94
rect -730 91 -726 94
rect -626 91 -622 94
rect -605 91 -601 94
rect -560 91 -556 94
rect -869 38 -865 41
rect -796 38 -792 41
rect -775 38 -771 41
rect -730 38 -726 41
rect -630 38 -626 41
rect -609 38 -605 41
rect -564 38 -560 41
rect -436 38 -432 41
rect -869 -1 -865 30
rect -796 -7 -792 30
rect -775 -7 -771 30
rect -730 -7 -726 30
rect -630 -7 -626 30
rect -609 -7 -605 30
rect -564 -7 -560 30
rect -869 -12 -865 -9
rect -436 -8 -432 30
rect -796 -18 -792 -15
rect -775 -18 -771 -15
rect -730 -18 -726 -15
rect -630 -18 -626 -15
rect -609 -18 -605 -15
rect -564 -18 -560 -15
rect -147 -16 -143 -13
rect -126 -16 -122 -13
rect 451 -16 455 -13
rect 472 -16 476 -13
rect 1330 -16 1334 -13
rect 1351 -16 1355 -13
rect 2098 -16 2102 -13
rect 2119 -16 2123 -13
rect -436 -19 -432 -16
rect -147 -61 -143 -24
rect -126 -61 -122 -24
rect 451 -61 455 -24
rect 472 -61 476 -24
rect 1330 -61 1334 -24
rect 1351 -61 1355 -24
rect 2098 -61 2102 -24
rect 2119 -61 2123 -24
rect -220 -64 -216 -61
rect -199 -64 -195 -61
rect 378 -64 382 -61
rect 399 -64 403 -61
rect -147 -72 -143 -69
rect -220 -109 -216 -72
rect -199 -109 -195 -72
rect -126 -76 -122 -69
rect 1257 -64 1261 -61
rect 1278 -64 1282 -61
rect 451 -72 455 -69
rect -46 -84 -42 -81
rect -25 -84 -21 -81
rect -574 -117 -570 -114
rect -553 -117 -549 -114
rect -508 -117 -504 -114
rect -220 -120 -216 -117
rect -199 -125 -195 -117
rect -132 -125 -128 -122
rect -111 -125 -107 -122
rect -574 -162 -570 -125
rect -553 -162 -549 -125
rect -508 -162 -504 -125
rect -46 -129 -42 -92
rect -25 -129 -21 -92
rect 378 -109 382 -72
rect 399 -109 403 -72
rect 472 -76 476 -69
rect 2025 -64 2029 -61
rect 2046 -64 2050 -61
rect 1330 -72 1334 -69
rect 552 -84 556 -81
rect 573 -84 577 -81
rect 378 -120 382 -117
rect 399 -125 403 -117
rect 466 -125 470 -122
rect 487 -125 491 -122
rect -132 -170 -128 -133
rect -111 -170 -107 -133
rect 552 -129 556 -92
rect 573 -129 577 -92
rect 1257 -109 1261 -72
rect 1278 -109 1282 -72
rect 1351 -76 1355 -69
rect 2098 -72 2102 -69
rect 1431 -84 1435 -81
rect 1452 -84 1456 -81
rect 1257 -120 1261 -117
rect 1278 -125 1282 -117
rect 1345 -125 1349 -122
rect 1366 -125 1370 -122
rect -46 -140 -42 -137
rect -25 -145 -21 -137
rect 466 -170 470 -133
rect 487 -170 491 -133
rect 1431 -129 1435 -92
rect 1452 -129 1456 -92
rect 2025 -109 2029 -72
rect 2046 -109 2050 -72
rect 2119 -76 2123 -69
rect 2199 -84 2203 -81
rect 2220 -84 2224 -81
rect 2025 -120 2029 -117
rect 2046 -125 2050 -117
rect 2113 -125 2117 -122
rect 2134 -125 2138 -122
rect 552 -140 556 -137
rect 573 -145 577 -137
rect 1345 -170 1349 -133
rect 1366 -170 1370 -133
rect 2199 -129 2203 -92
rect 2220 -129 2224 -92
rect 1431 -140 1435 -137
rect 1452 -145 1456 -137
rect 2113 -170 2117 -133
rect 2134 -170 2138 -133
rect 2199 -140 2203 -137
rect 2220 -145 2224 -137
rect -574 -173 -570 -170
rect -553 -173 -549 -170
rect -508 -173 -504 -170
rect -132 -181 -128 -178
rect -111 -186 -107 -178
rect 466 -181 470 -178
rect 487 -186 491 -178
rect 1345 -181 1349 -178
rect 1366 -186 1370 -178
rect 2113 -181 2117 -178
rect 2134 -186 2138 -178
rect -577 -209 -573 -206
rect -556 -209 -552 -206
rect -511 -209 -507 -206
rect -577 -254 -573 -217
rect -556 -254 -552 -217
rect -511 -254 -507 -217
rect -577 -265 -573 -262
rect -556 -265 -552 -262
rect -511 -265 -507 -262
rect -577 -301 -573 -298
rect -556 -301 -552 -298
rect -511 -301 -507 -298
rect -577 -346 -573 -309
rect -556 -346 -552 -309
rect -511 -346 -507 -309
rect 134 -319 138 -316
rect 155 -319 159 -316
rect 877 -322 881 -319
rect 898 -322 902 -319
rect 1636 -322 1640 -319
rect 1657 -322 1661 -319
rect 2372 -322 2376 -319
rect 2393 -322 2397 -319
rect -577 -357 -573 -354
rect -556 -357 -552 -354
rect -511 -357 -507 -354
rect 134 -364 138 -327
rect 155 -364 159 -327
rect -176 -367 -172 -364
rect -155 -367 -151 -364
rect 61 -367 65 -364
rect 82 -367 86 -364
rect 877 -367 881 -330
rect 898 -367 902 -330
rect 1636 -367 1640 -330
rect 1657 -367 1661 -330
rect 2372 -367 2376 -330
rect 2393 -367 2397 -330
rect 567 -370 571 -367
rect 588 -370 592 -367
rect 804 -370 808 -367
rect 825 -370 829 -367
rect 134 -375 138 -372
rect -577 -393 -573 -390
rect -556 -393 -552 -390
rect -511 -393 -507 -390
rect -577 -438 -573 -401
rect -556 -438 -552 -401
rect -511 -438 -507 -401
rect -176 -412 -172 -375
rect -155 -412 -151 -375
rect 61 -412 65 -375
rect 82 -412 86 -375
rect 155 -379 159 -372
rect 1326 -370 1330 -367
rect 1347 -370 1351 -367
rect 1563 -370 1567 -367
rect 1584 -370 1588 -367
rect 877 -378 881 -375
rect 235 -387 239 -384
rect 256 -387 260 -384
rect -249 -415 -245 -412
rect -228 -415 -224 -412
rect -176 -423 -172 -420
rect -577 -449 -573 -446
rect -556 -449 -552 -446
rect -511 -449 -507 -446
rect -249 -460 -245 -423
rect -228 -460 -224 -423
rect -155 -427 -151 -420
rect 61 -423 65 -420
rect 82 -428 86 -420
rect 149 -428 153 -425
rect 170 -428 174 -425
rect -75 -435 -71 -432
rect -54 -435 -50 -432
rect 235 -432 239 -395
rect 256 -432 260 -395
rect 567 -415 571 -378
rect 588 -415 592 -378
rect 804 -415 808 -378
rect 825 -415 829 -378
rect 898 -382 902 -375
rect 2062 -370 2066 -367
rect 2083 -370 2087 -367
rect 2299 -370 2303 -367
rect 2320 -370 2324 -367
rect 1636 -378 1640 -375
rect 978 -390 982 -387
rect 999 -390 1003 -387
rect 494 -418 498 -415
rect 515 -418 519 -415
rect 567 -426 571 -423
rect -249 -471 -245 -468
rect -228 -476 -224 -468
rect -161 -476 -157 -473
rect -140 -476 -136 -473
rect -572 -484 -568 -481
rect -551 -484 -547 -481
rect -506 -484 -502 -481
rect -75 -480 -71 -443
rect -54 -480 -50 -443
rect 149 -473 153 -436
rect 170 -473 174 -436
rect 235 -443 239 -440
rect 256 -448 260 -440
rect 494 -463 498 -426
rect 515 -463 519 -426
rect 588 -430 592 -423
rect 804 -426 808 -423
rect 825 -431 829 -423
rect 892 -431 896 -428
rect 913 -431 917 -428
rect 668 -438 672 -435
rect 689 -438 693 -435
rect 978 -435 982 -398
rect 999 -435 1003 -398
rect 1326 -415 1330 -378
rect 1347 -415 1351 -378
rect 1563 -415 1567 -378
rect 1584 -415 1588 -378
rect 1657 -382 1661 -375
rect 2372 -378 2376 -375
rect 1737 -390 1741 -387
rect 1758 -390 1762 -387
rect 1253 -418 1257 -415
rect 1274 -418 1278 -415
rect 1326 -426 1330 -423
rect -572 -529 -568 -492
rect -551 -529 -547 -492
rect -506 -529 -502 -492
rect -161 -521 -157 -484
rect -140 -521 -136 -484
rect 494 -474 498 -471
rect 515 -479 519 -471
rect 582 -479 586 -476
rect 603 -479 607 -476
rect 149 -484 153 -481
rect -75 -491 -71 -488
rect -54 -496 -50 -488
rect 170 -489 174 -481
rect 668 -483 672 -446
rect 689 -483 693 -446
rect 892 -476 896 -439
rect 913 -476 917 -439
rect 978 -446 982 -443
rect 999 -451 1003 -443
rect 1253 -463 1257 -426
rect 1274 -463 1278 -426
rect 1347 -430 1351 -423
rect 1563 -426 1567 -423
rect 1584 -431 1588 -423
rect 1651 -431 1655 -428
rect 1672 -431 1676 -428
rect 1427 -438 1431 -435
rect 1448 -438 1452 -435
rect 1737 -435 1741 -398
rect 1758 -435 1762 -398
rect 2062 -415 2066 -378
rect 2083 -415 2087 -378
rect 2299 -415 2303 -378
rect 2320 -415 2324 -378
rect 2393 -382 2397 -375
rect 2473 -390 2477 -387
rect 2494 -390 2498 -387
rect 1989 -418 1993 -415
rect 2010 -418 2014 -415
rect 2062 -426 2066 -423
rect 1253 -474 1257 -471
rect 582 -524 586 -487
rect 603 -524 607 -487
rect 1274 -479 1278 -471
rect 1341 -479 1345 -476
rect 1362 -479 1366 -476
rect 892 -487 896 -484
rect 668 -494 672 -491
rect 689 -499 693 -491
rect 913 -492 917 -484
rect 1427 -483 1431 -446
rect 1448 -483 1452 -446
rect 1651 -476 1655 -439
rect 1672 -476 1676 -439
rect 1737 -446 1741 -443
rect 1758 -451 1762 -443
rect 1989 -463 1993 -426
rect 2010 -463 2014 -426
rect 2083 -430 2087 -423
rect 2299 -426 2303 -423
rect 2320 -431 2324 -423
rect 2387 -431 2391 -428
rect 2408 -431 2412 -428
rect 2163 -438 2167 -435
rect 2184 -438 2188 -435
rect 2473 -435 2477 -398
rect 2494 -435 2498 -398
rect 1989 -474 1993 -471
rect 1341 -524 1345 -487
rect 1362 -524 1366 -487
rect 2010 -479 2014 -471
rect 2077 -479 2081 -476
rect 2098 -479 2102 -476
rect 1651 -487 1655 -484
rect 1427 -494 1431 -491
rect 1448 -499 1452 -491
rect 1672 -492 1676 -484
rect 2163 -483 2167 -446
rect 2184 -483 2188 -446
rect 2387 -476 2391 -439
rect 2408 -476 2412 -439
rect 2473 -446 2477 -443
rect 2494 -451 2498 -443
rect 2077 -524 2081 -487
rect 2098 -524 2102 -487
rect 2387 -487 2391 -484
rect 2163 -494 2167 -491
rect 2184 -499 2188 -491
rect 2408 -492 2412 -484
rect -161 -532 -157 -529
rect -140 -537 -136 -529
rect 121 -534 125 -531
rect 142 -534 146 -531
rect 187 -534 191 -531
rect 280 -534 284 -531
rect 301 -534 305 -531
rect 348 -534 352 -531
rect -572 -540 -568 -537
rect -551 -540 -547 -537
rect -506 -540 -502 -537
rect 582 -535 586 -532
rect 603 -540 607 -532
rect 864 -537 868 -534
rect 885 -537 889 -534
rect 930 -537 934 -534
rect 1023 -537 1027 -534
rect 1044 -537 1048 -534
rect 1091 -537 1095 -534
rect 1341 -535 1345 -532
rect -575 -576 -571 -573
rect -554 -576 -550 -573
rect -509 -576 -505 -573
rect 121 -579 125 -542
rect 142 -579 146 -542
rect 187 -579 191 -542
rect -575 -621 -571 -584
rect -554 -621 -550 -584
rect -509 -621 -505 -584
rect -190 -585 -186 -582
rect -169 -585 -165 -582
rect -124 -585 -120 -582
rect 280 -582 284 -542
rect 301 -582 305 -542
rect 348 -582 352 -542
rect 1362 -540 1366 -532
rect 1623 -537 1627 -534
rect 1644 -537 1648 -534
rect 1689 -537 1693 -534
rect 1782 -537 1786 -534
rect 1803 -537 1807 -534
rect 1850 -537 1854 -534
rect 2077 -535 2081 -532
rect 2098 -540 2102 -532
rect 2359 -537 2363 -534
rect 2380 -537 2384 -534
rect 2425 -537 2429 -534
rect 2518 -537 2522 -534
rect 2539 -537 2543 -534
rect 2586 -537 2590 -534
rect 864 -582 868 -545
rect 885 -582 889 -545
rect 930 -582 934 -545
rect 121 -590 125 -587
rect 142 -590 146 -587
rect 187 -590 191 -587
rect 553 -588 557 -585
rect 574 -588 578 -585
rect 619 -588 623 -585
rect 280 -593 284 -590
rect 301 -593 305 -590
rect 348 -593 352 -590
rect -575 -632 -571 -629
rect -554 -632 -550 -629
rect -509 -632 -505 -629
rect -190 -630 -186 -593
rect -169 -630 -165 -593
rect -124 -630 -120 -593
rect 1023 -585 1027 -545
rect 1044 -585 1048 -545
rect 1091 -585 1095 -545
rect 1623 -582 1627 -545
rect 1644 -582 1648 -545
rect 1689 -582 1693 -545
rect 864 -593 868 -590
rect 885 -593 889 -590
rect 930 -593 934 -590
rect 1312 -588 1316 -585
rect 1333 -588 1337 -585
rect 1378 -588 1382 -585
rect 1023 -596 1027 -593
rect 1044 -596 1048 -593
rect 1091 -596 1095 -593
rect 1782 -585 1786 -545
rect 1803 -585 1807 -545
rect 1850 -585 1854 -545
rect 2359 -582 2363 -545
rect 2380 -582 2384 -545
rect 2425 -582 2429 -545
rect 1623 -593 1627 -590
rect 1644 -593 1648 -590
rect 1689 -593 1693 -590
rect 2048 -588 2052 -585
rect 2069 -588 2073 -585
rect 2114 -588 2118 -585
rect 1782 -596 1786 -593
rect 1803 -596 1807 -593
rect 1850 -596 1854 -593
rect 2518 -585 2522 -545
rect 2539 -585 2543 -545
rect 2586 -585 2590 -545
rect 2359 -593 2363 -590
rect 2380 -593 2384 -590
rect 2425 -593 2429 -590
rect 2518 -596 2522 -593
rect 2539 -596 2543 -593
rect 2586 -596 2590 -593
rect 553 -633 557 -596
rect 574 -633 578 -596
rect 619 -633 623 -596
rect 1312 -633 1316 -596
rect 1333 -633 1337 -596
rect 1378 -633 1382 -596
rect 2048 -633 2052 -596
rect 2069 -633 2073 -596
rect 2114 -633 2118 -596
rect -190 -641 -186 -638
rect -169 -641 -165 -638
rect -124 -641 -120 -638
rect 553 -644 557 -641
rect 574 -644 578 -641
rect 619 -644 623 -641
rect 1312 -644 1316 -641
rect 1333 -644 1337 -641
rect 1378 -644 1382 -641
rect 2048 -644 2052 -641
rect 2069 -644 2073 -641
rect 2114 -644 2118 -641
rect -575 -668 -571 -665
rect -554 -668 -550 -665
rect -509 -668 -505 -665
rect -575 -713 -571 -676
rect -554 -713 -550 -676
rect -509 -713 -505 -676
rect -575 -724 -571 -721
rect -554 -724 -550 -721
rect -509 -724 -505 -721
rect -575 -760 -571 -757
rect -554 -760 -550 -757
rect -509 -760 -505 -757
rect -575 -805 -571 -768
rect -554 -805 -550 -768
rect -509 -805 -505 -768
rect -118 -809 -114 -806
rect -97 -809 -93 -806
rect 480 -809 484 -806
rect 501 -809 505 -806
rect 1359 -809 1363 -806
rect 1380 -809 1384 -806
rect 2127 -809 2131 -806
rect 2148 -809 2152 -806
rect -575 -816 -571 -813
rect -554 -816 -550 -813
rect -509 -816 -505 -813
rect -118 -854 -114 -817
rect -97 -854 -93 -817
rect 480 -854 484 -817
rect 501 -854 505 -817
rect 1359 -854 1363 -817
rect 1380 -854 1384 -817
rect 2127 -854 2131 -817
rect 2148 -854 2152 -817
rect -191 -857 -187 -854
rect -170 -857 -166 -854
rect 407 -857 411 -854
rect 428 -857 432 -854
rect -118 -865 -114 -862
rect -191 -902 -187 -865
rect -170 -902 -166 -865
rect -97 -869 -93 -862
rect 1286 -857 1290 -854
rect 1307 -857 1311 -854
rect 480 -865 484 -862
rect -17 -877 -13 -874
rect 4 -877 8 -874
rect -574 -910 -570 -907
rect -553 -910 -549 -907
rect -508 -910 -504 -907
rect -191 -913 -187 -910
rect -170 -918 -166 -910
rect -103 -918 -99 -915
rect -82 -918 -78 -915
rect -574 -955 -570 -918
rect -553 -955 -549 -918
rect -508 -955 -504 -918
rect -17 -922 -13 -885
rect 4 -922 8 -885
rect 407 -902 411 -865
rect 428 -902 432 -865
rect 501 -869 505 -862
rect 2054 -857 2058 -854
rect 2075 -857 2079 -854
rect 1359 -865 1363 -862
rect 581 -877 585 -874
rect 602 -877 606 -874
rect 407 -913 411 -910
rect 428 -918 432 -910
rect 495 -918 499 -915
rect 516 -918 520 -915
rect -103 -963 -99 -926
rect -82 -963 -78 -926
rect 581 -922 585 -885
rect 602 -922 606 -885
rect 1286 -902 1290 -865
rect 1307 -902 1311 -865
rect 1380 -869 1384 -862
rect 2127 -865 2131 -862
rect 1460 -877 1464 -874
rect 1481 -877 1485 -874
rect 1286 -913 1290 -910
rect 1307 -918 1311 -910
rect 1374 -918 1378 -915
rect 1395 -918 1399 -915
rect -17 -933 -13 -930
rect 4 -938 8 -930
rect 495 -963 499 -926
rect 516 -963 520 -926
rect 1460 -922 1464 -885
rect 1481 -922 1485 -885
rect 2054 -902 2058 -865
rect 2075 -902 2079 -865
rect 2148 -869 2152 -862
rect 2228 -877 2232 -874
rect 2249 -877 2253 -874
rect 2054 -913 2058 -910
rect 2075 -918 2079 -910
rect 2142 -918 2146 -915
rect 2163 -918 2167 -915
rect 581 -933 585 -930
rect 602 -938 606 -930
rect 1374 -963 1378 -926
rect 1395 -963 1399 -926
rect 2228 -922 2232 -885
rect 2249 -922 2253 -885
rect 1460 -933 1464 -930
rect 1481 -938 1485 -930
rect 2142 -963 2146 -926
rect 2163 -963 2167 -926
rect 2228 -933 2232 -930
rect 2249 -938 2253 -930
rect -574 -966 -570 -963
rect -553 -966 -549 -963
rect -508 -966 -504 -963
rect -103 -974 -99 -971
rect -82 -979 -78 -971
rect 495 -974 499 -971
rect 516 -979 520 -971
rect 1374 -974 1378 -971
rect 1395 -979 1399 -971
rect 2142 -974 2146 -971
rect 2163 -979 2167 -971
rect -577 -1002 -573 -999
rect -556 -1002 -552 -999
rect -511 -1002 -507 -999
rect -577 -1047 -573 -1010
rect -556 -1047 -552 -1010
rect -511 -1047 -507 -1010
rect -577 -1058 -573 -1055
rect -556 -1058 -552 -1055
rect -511 -1058 -507 -1055
rect -577 -1094 -573 -1091
rect -556 -1094 -552 -1091
rect -511 -1094 -507 -1091
rect -577 -1139 -573 -1102
rect -556 -1139 -552 -1102
rect -511 -1139 -507 -1102
rect 163 -1112 167 -1109
rect 184 -1112 188 -1109
rect 906 -1115 910 -1112
rect 927 -1115 931 -1112
rect 1665 -1115 1669 -1112
rect 1686 -1115 1690 -1112
rect 2401 -1115 2405 -1112
rect 2422 -1115 2426 -1112
rect -577 -1150 -573 -1147
rect -556 -1150 -552 -1147
rect -511 -1150 -507 -1147
rect 163 -1157 167 -1120
rect 184 -1157 188 -1120
rect -147 -1160 -143 -1157
rect -126 -1160 -122 -1157
rect 90 -1160 94 -1157
rect 111 -1160 115 -1157
rect 906 -1160 910 -1123
rect 927 -1160 931 -1123
rect 1665 -1160 1669 -1123
rect 1686 -1160 1690 -1123
rect 2401 -1160 2405 -1123
rect 2422 -1160 2426 -1123
rect 596 -1163 600 -1160
rect 617 -1163 621 -1160
rect 833 -1163 837 -1160
rect 854 -1163 858 -1160
rect 163 -1168 167 -1165
rect -577 -1186 -573 -1183
rect -556 -1186 -552 -1183
rect -511 -1186 -507 -1183
rect -577 -1231 -573 -1194
rect -556 -1231 -552 -1194
rect -511 -1231 -507 -1194
rect -147 -1205 -143 -1168
rect -126 -1205 -122 -1168
rect 90 -1205 94 -1168
rect 111 -1205 115 -1168
rect 184 -1172 188 -1165
rect 1355 -1163 1359 -1160
rect 1376 -1163 1380 -1160
rect 1592 -1163 1596 -1160
rect 1613 -1163 1617 -1160
rect 906 -1171 910 -1168
rect 264 -1180 268 -1177
rect 285 -1180 289 -1177
rect -220 -1208 -216 -1205
rect -199 -1208 -195 -1205
rect -147 -1216 -143 -1213
rect -577 -1242 -573 -1239
rect -556 -1242 -552 -1239
rect -511 -1242 -507 -1239
rect -220 -1253 -216 -1216
rect -199 -1253 -195 -1216
rect -126 -1220 -122 -1213
rect 90 -1216 94 -1213
rect 111 -1221 115 -1213
rect 178 -1221 182 -1218
rect 199 -1221 203 -1218
rect -46 -1228 -42 -1225
rect -25 -1228 -21 -1225
rect 264 -1225 268 -1188
rect 285 -1225 289 -1188
rect 596 -1208 600 -1171
rect 617 -1208 621 -1171
rect 833 -1208 837 -1171
rect 854 -1208 858 -1171
rect 927 -1175 931 -1168
rect 2091 -1163 2095 -1160
rect 2112 -1163 2116 -1160
rect 2328 -1163 2332 -1160
rect 2349 -1163 2353 -1160
rect 1665 -1171 1669 -1168
rect 1007 -1183 1011 -1180
rect 1028 -1183 1032 -1180
rect 523 -1211 527 -1208
rect 544 -1211 548 -1208
rect 596 -1219 600 -1216
rect -220 -1264 -216 -1261
rect -199 -1269 -195 -1261
rect -132 -1269 -128 -1266
rect -111 -1269 -107 -1266
rect -572 -1277 -568 -1274
rect -551 -1277 -547 -1274
rect -506 -1277 -502 -1274
rect -46 -1273 -42 -1236
rect -25 -1273 -21 -1236
rect 178 -1266 182 -1229
rect 199 -1266 203 -1229
rect 264 -1236 268 -1233
rect 285 -1241 289 -1233
rect 523 -1256 527 -1219
rect 544 -1256 548 -1219
rect 617 -1223 621 -1216
rect 833 -1219 837 -1216
rect 854 -1224 858 -1216
rect 921 -1224 925 -1221
rect 942 -1224 946 -1221
rect 697 -1231 701 -1228
rect 718 -1231 722 -1228
rect 1007 -1228 1011 -1191
rect 1028 -1228 1032 -1191
rect 1355 -1208 1359 -1171
rect 1376 -1208 1380 -1171
rect 1592 -1208 1596 -1171
rect 1613 -1208 1617 -1171
rect 1686 -1175 1690 -1168
rect 2401 -1171 2405 -1168
rect 1766 -1183 1770 -1180
rect 1787 -1183 1791 -1180
rect 1282 -1211 1286 -1208
rect 1303 -1211 1307 -1208
rect 1355 -1219 1359 -1216
rect -572 -1322 -568 -1285
rect -551 -1322 -547 -1285
rect -506 -1322 -502 -1285
rect -132 -1314 -128 -1277
rect -111 -1314 -107 -1277
rect 523 -1267 527 -1264
rect 544 -1272 548 -1264
rect 611 -1272 615 -1269
rect 632 -1272 636 -1269
rect 178 -1277 182 -1274
rect -46 -1284 -42 -1281
rect -25 -1289 -21 -1281
rect 199 -1282 203 -1274
rect 697 -1276 701 -1239
rect 718 -1276 722 -1239
rect 921 -1269 925 -1232
rect 942 -1269 946 -1232
rect 1007 -1239 1011 -1236
rect 1028 -1244 1032 -1236
rect 1282 -1256 1286 -1219
rect 1303 -1256 1307 -1219
rect 1376 -1223 1380 -1216
rect 1592 -1219 1596 -1216
rect 1613 -1224 1617 -1216
rect 1680 -1224 1684 -1221
rect 1701 -1224 1705 -1221
rect 1456 -1231 1460 -1228
rect 1477 -1231 1481 -1228
rect 1766 -1228 1770 -1191
rect 1787 -1228 1791 -1191
rect 2091 -1208 2095 -1171
rect 2112 -1208 2116 -1171
rect 2328 -1208 2332 -1171
rect 2349 -1208 2353 -1171
rect 2422 -1175 2426 -1168
rect 2502 -1183 2506 -1180
rect 2523 -1183 2527 -1180
rect 2018 -1211 2022 -1208
rect 2039 -1211 2043 -1208
rect 2091 -1219 2095 -1216
rect 1282 -1267 1286 -1264
rect 611 -1317 615 -1280
rect 632 -1317 636 -1280
rect 1303 -1272 1307 -1264
rect 1370 -1272 1374 -1269
rect 1391 -1272 1395 -1269
rect 921 -1280 925 -1277
rect 697 -1287 701 -1284
rect 718 -1292 722 -1284
rect 942 -1285 946 -1277
rect 1456 -1276 1460 -1239
rect 1477 -1276 1481 -1239
rect 1680 -1269 1684 -1232
rect 1701 -1269 1705 -1232
rect 1766 -1239 1770 -1236
rect 1787 -1244 1791 -1236
rect 2018 -1256 2022 -1219
rect 2039 -1256 2043 -1219
rect 2112 -1223 2116 -1216
rect 2328 -1219 2332 -1216
rect 2349 -1224 2353 -1216
rect 2416 -1224 2420 -1221
rect 2437 -1224 2441 -1221
rect 2192 -1231 2196 -1228
rect 2213 -1231 2217 -1228
rect 2502 -1228 2506 -1191
rect 2523 -1228 2527 -1191
rect 2018 -1267 2022 -1264
rect 1370 -1317 1374 -1280
rect 1391 -1317 1395 -1280
rect 2039 -1272 2043 -1264
rect 2106 -1272 2110 -1269
rect 2127 -1272 2131 -1269
rect 1680 -1280 1684 -1277
rect 1456 -1287 1460 -1284
rect 1477 -1292 1481 -1284
rect 1701 -1285 1705 -1277
rect 2192 -1276 2196 -1239
rect 2213 -1276 2217 -1239
rect 2416 -1269 2420 -1232
rect 2437 -1269 2441 -1232
rect 2502 -1239 2506 -1236
rect 2523 -1244 2527 -1236
rect 2106 -1317 2110 -1280
rect 2127 -1317 2131 -1280
rect 2416 -1280 2420 -1277
rect 2192 -1287 2196 -1284
rect 2213 -1292 2217 -1284
rect 2437 -1285 2441 -1277
rect -132 -1325 -128 -1322
rect -111 -1330 -107 -1322
rect 150 -1327 154 -1324
rect 171 -1327 175 -1324
rect 216 -1327 220 -1324
rect 309 -1327 313 -1324
rect 330 -1327 334 -1324
rect 377 -1327 381 -1324
rect -572 -1333 -568 -1330
rect -551 -1333 -547 -1330
rect -506 -1333 -502 -1330
rect 611 -1328 615 -1325
rect 632 -1333 636 -1325
rect 893 -1330 897 -1327
rect 914 -1330 918 -1327
rect 959 -1330 963 -1327
rect 1052 -1330 1056 -1327
rect 1073 -1330 1077 -1327
rect 1120 -1330 1124 -1327
rect 1370 -1328 1374 -1325
rect -575 -1369 -571 -1366
rect -554 -1369 -550 -1366
rect -509 -1369 -505 -1366
rect 150 -1372 154 -1335
rect 171 -1372 175 -1335
rect 216 -1372 220 -1335
rect -575 -1414 -571 -1377
rect -554 -1414 -550 -1377
rect -509 -1414 -505 -1377
rect -161 -1378 -157 -1375
rect -140 -1378 -136 -1375
rect -95 -1378 -91 -1375
rect 309 -1375 313 -1335
rect 330 -1375 334 -1335
rect 377 -1375 381 -1335
rect 1391 -1333 1395 -1325
rect 1652 -1330 1656 -1327
rect 1673 -1330 1677 -1327
rect 1718 -1330 1722 -1327
rect 1811 -1330 1815 -1327
rect 1832 -1330 1836 -1327
rect 1879 -1330 1883 -1327
rect 2106 -1328 2110 -1325
rect 2127 -1333 2131 -1325
rect 2388 -1330 2392 -1327
rect 2409 -1330 2413 -1327
rect 2454 -1330 2458 -1327
rect 2547 -1330 2551 -1327
rect 2568 -1330 2572 -1327
rect 2615 -1330 2619 -1327
rect 893 -1375 897 -1338
rect 914 -1375 918 -1338
rect 959 -1375 963 -1338
rect 150 -1383 154 -1380
rect 171 -1383 175 -1380
rect 216 -1383 220 -1380
rect 582 -1381 586 -1378
rect 603 -1381 607 -1378
rect 648 -1381 652 -1378
rect 309 -1386 313 -1383
rect 330 -1386 334 -1383
rect 377 -1386 381 -1383
rect -575 -1425 -571 -1422
rect -554 -1425 -550 -1422
rect -509 -1425 -505 -1422
rect -161 -1423 -157 -1386
rect -140 -1423 -136 -1386
rect -95 -1423 -91 -1386
rect 1052 -1378 1056 -1338
rect 1073 -1378 1077 -1338
rect 1120 -1378 1124 -1338
rect 1652 -1375 1656 -1338
rect 1673 -1375 1677 -1338
rect 1718 -1375 1722 -1338
rect 893 -1386 897 -1383
rect 914 -1386 918 -1383
rect 959 -1386 963 -1383
rect 1341 -1381 1345 -1378
rect 1362 -1381 1366 -1378
rect 1407 -1381 1411 -1378
rect 1052 -1389 1056 -1386
rect 1073 -1389 1077 -1386
rect 1120 -1389 1124 -1386
rect 1811 -1378 1815 -1338
rect 1832 -1378 1836 -1338
rect 1879 -1378 1883 -1338
rect 2388 -1375 2392 -1338
rect 2409 -1375 2413 -1338
rect 2454 -1375 2458 -1338
rect 1652 -1386 1656 -1383
rect 1673 -1386 1677 -1383
rect 1718 -1386 1722 -1383
rect 2077 -1381 2081 -1378
rect 2098 -1381 2102 -1378
rect 2143 -1381 2147 -1378
rect 1811 -1389 1815 -1386
rect 1832 -1389 1836 -1386
rect 1879 -1389 1883 -1386
rect 2547 -1378 2551 -1338
rect 2568 -1378 2572 -1338
rect 2615 -1378 2619 -1338
rect 2388 -1386 2392 -1383
rect 2409 -1386 2413 -1383
rect 2454 -1386 2458 -1383
rect 2547 -1389 2551 -1386
rect 2568 -1389 2572 -1386
rect 2615 -1389 2619 -1386
rect 582 -1426 586 -1389
rect 603 -1426 607 -1389
rect 648 -1426 652 -1389
rect 1341 -1426 1345 -1389
rect 1362 -1426 1366 -1389
rect 1407 -1426 1411 -1389
rect 2077 -1426 2081 -1389
rect 2098 -1426 2102 -1389
rect 2143 -1426 2147 -1389
rect -161 -1434 -157 -1431
rect -140 -1434 -136 -1431
rect -95 -1434 -91 -1431
rect 582 -1437 586 -1434
rect 603 -1437 607 -1434
rect 648 -1437 652 -1434
rect 1341 -1437 1345 -1434
rect 1362 -1437 1366 -1434
rect 1407 -1437 1411 -1434
rect 2077 -1437 2081 -1434
rect 2098 -1437 2102 -1434
rect 2143 -1437 2147 -1434
rect -575 -1461 -571 -1458
rect -554 -1461 -550 -1458
rect -509 -1461 -505 -1458
rect -575 -1506 -571 -1469
rect -554 -1506 -550 -1469
rect -509 -1506 -505 -1469
rect -575 -1517 -571 -1514
rect -554 -1517 -550 -1514
rect -509 -1517 -505 -1514
rect -575 -1553 -571 -1550
rect -554 -1553 -550 -1550
rect -509 -1553 -505 -1550
rect -575 -1598 -571 -1561
rect -554 -1598 -550 -1561
rect -509 -1598 -505 -1561
rect -575 -1609 -571 -1606
rect -554 -1609 -550 -1606
rect -509 -1609 -505 -1606
rect -574 -1673 -570 -1670
rect -553 -1673 -549 -1670
rect -508 -1673 -504 -1670
rect -574 -1718 -570 -1681
rect -553 -1718 -549 -1681
rect -508 -1718 -504 -1681
rect -574 -1729 -570 -1726
rect -553 -1729 -549 -1726
rect -508 -1729 -504 -1726
rect 19 -1729 23 -1726
rect 40 -1729 44 -1726
rect 508 -1729 512 -1726
rect 529 -1729 533 -1726
rect 892 -1729 896 -1726
rect 913 -1729 917 -1726
rect -577 -1765 -573 -1762
rect -556 -1765 -552 -1762
rect -511 -1765 -507 -1762
rect -577 -1810 -573 -1773
rect -556 -1810 -552 -1773
rect -511 -1810 -507 -1773
rect 19 -1774 23 -1737
rect 40 -1774 44 -1737
rect 508 -1774 512 -1737
rect 529 -1774 533 -1737
rect 892 -1774 896 -1737
rect 913 -1774 917 -1737
rect 1307 -1753 1311 -1750
rect 1328 -1753 1332 -1750
rect -54 -1777 -50 -1774
rect -33 -1777 -29 -1774
rect 435 -1777 439 -1774
rect 456 -1777 460 -1774
rect 19 -1785 23 -1782
rect -577 -1821 -573 -1818
rect -556 -1821 -552 -1818
rect -511 -1821 -507 -1818
rect -54 -1822 -50 -1785
rect -33 -1822 -29 -1785
rect 40 -1789 44 -1782
rect 819 -1777 823 -1774
rect 840 -1777 844 -1774
rect 508 -1785 512 -1782
rect 120 -1797 124 -1794
rect 141 -1797 145 -1794
rect 246 -1801 250 -1798
rect -54 -1833 -50 -1830
rect -33 -1838 -29 -1830
rect 34 -1838 38 -1835
rect 55 -1838 59 -1835
rect 120 -1842 124 -1805
rect 141 -1842 145 -1805
rect 246 -1840 250 -1809
rect 435 -1822 439 -1785
rect 456 -1822 460 -1785
rect 529 -1789 533 -1782
rect 892 -1785 896 -1782
rect 609 -1797 613 -1794
rect 630 -1797 634 -1794
rect 682 -1801 686 -1798
rect 435 -1833 439 -1830
rect 456 -1838 460 -1830
rect 523 -1838 527 -1835
rect 544 -1838 548 -1835
rect -577 -1857 -573 -1854
rect -556 -1857 -552 -1854
rect -511 -1857 -507 -1854
rect -577 -1902 -573 -1865
rect -556 -1902 -552 -1865
rect -511 -1902 -507 -1865
rect 34 -1883 38 -1846
rect 55 -1883 59 -1846
rect 609 -1842 613 -1805
rect 630 -1842 634 -1805
rect 682 -1840 686 -1809
rect 819 -1822 823 -1785
rect 840 -1822 844 -1785
rect 913 -1789 917 -1782
rect 1027 -1797 1031 -1794
rect 1048 -1797 1052 -1794
rect 1307 -1798 1311 -1761
rect 1328 -1798 1332 -1761
rect 1100 -1801 1104 -1798
rect 1234 -1801 1238 -1798
rect 1255 -1801 1259 -1798
rect 819 -1833 823 -1830
rect 840 -1838 844 -1830
rect 907 -1838 911 -1835
rect 928 -1838 932 -1835
rect 120 -1853 124 -1850
rect 141 -1858 145 -1850
rect 246 -1851 250 -1848
rect 523 -1883 527 -1846
rect 544 -1883 548 -1846
rect 1027 -1842 1031 -1805
rect 1048 -1842 1052 -1805
rect 1307 -1809 1311 -1806
rect 1100 -1840 1104 -1809
rect 609 -1853 613 -1850
rect 630 -1858 634 -1850
rect 682 -1851 686 -1848
rect 907 -1883 911 -1846
rect 928 -1883 932 -1846
rect 1234 -1846 1238 -1809
rect 1255 -1846 1259 -1809
rect 1328 -1813 1332 -1806
rect 1408 -1821 1412 -1818
rect 1429 -1821 1433 -1818
rect 1476 -1821 1480 -1818
rect 1027 -1853 1031 -1850
rect 1048 -1858 1052 -1850
rect 1100 -1851 1104 -1848
rect 1234 -1857 1238 -1854
rect 1255 -1862 1259 -1854
rect 1322 -1862 1326 -1859
rect 1343 -1862 1347 -1859
rect 1408 -1866 1412 -1829
rect 1429 -1866 1433 -1829
rect 1476 -1860 1480 -1829
rect 34 -1894 38 -1891
rect 55 -1899 59 -1891
rect 523 -1894 527 -1891
rect 544 -1899 548 -1891
rect 907 -1894 911 -1891
rect 928 -1899 932 -1891
rect 1322 -1907 1326 -1870
rect 1343 -1907 1347 -1870
rect 1476 -1871 1480 -1868
rect 1408 -1877 1412 -1874
rect 1429 -1882 1433 -1874
rect -577 -1913 -573 -1910
rect -556 -1913 -552 -1910
rect -511 -1913 -507 -1910
rect 1322 -1918 1326 -1915
rect 1343 -1923 1347 -1915
rect -577 -1949 -573 -1946
rect -556 -1949 -552 -1946
rect -511 -1949 -507 -1946
rect -577 -1994 -573 -1957
rect -556 -1994 -552 -1957
rect -511 -1994 -507 -1957
rect -577 -2005 -573 -2002
rect -556 -2005 -552 -2002
rect -511 -2005 -507 -2002
rect -572 -2040 -568 -2037
rect -551 -2040 -547 -2037
rect -506 -2040 -502 -2037
rect -572 -2085 -568 -2048
rect -551 -2085 -547 -2048
rect -506 -2085 -502 -2048
rect 339 -2087 343 -2084
rect 372 -2087 376 -2084
rect 396 -2087 400 -2084
rect 447 -2087 451 -2084
rect 755 -2087 759 -2084
rect 788 -2087 792 -2084
rect 812 -2087 816 -2084
rect 863 -2087 867 -2084
rect 1205 -2087 1209 -2084
rect 1238 -2087 1242 -2084
rect 1262 -2087 1266 -2084
rect 1313 -2087 1317 -2084
rect -572 -2096 -568 -2093
rect -551 -2096 -547 -2093
rect -506 -2096 -502 -2093
rect -575 -2132 -571 -2129
rect -554 -2132 -550 -2129
rect -509 -2132 -505 -2129
rect 261 -2140 265 -2137
rect -575 -2177 -571 -2140
rect -554 -2177 -550 -2140
rect -509 -2177 -505 -2140
rect -28 -2164 -24 -2161
rect 59 -2172 63 -2169
rect 80 -2172 84 -2169
rect 125 -2172 129 -2169
rect -575 -2188 -571 -2185
rect -554 -2188 -550 -2185
rect -509 -2188 -505 -2185
rect -28 -2203 -24 -2172
rect -28 -2214 -24 -2211
rect 59 -2217 63 -2180
rect 80 -2217 84 -2180
rect 125 -2217 129 -2180
rect 261 -2185 265 -2148
rect 339 -2161 343 -2095
rect 372 -2161 376 -2095
rect 396 -2161 400 -2095
rect 447 -2161 451 -2095
rect 677 -2140 681 -2137
rect 339 -2172 343 -2169
rect 372 -2172 376 -2169
rect 396 -2172 400 -2169
rect 447 -2172 451 -2169
rect 677 -2185 681 -2148
rect 755 -2161 759 -2095
rect 788 -2161 792 -2095
rect 812 -2161 816 -2095
rect 863 -2161 867 -2095
rect 1121 -2140 1125 -2137
rect 755 -2172 759 -2169
rect 788 -2172 792 -2169
rect 812 -2172 816 -2169
rect 863 -2172 867 -2169
rect 1121 -2185 1125 -2148
rect 1205 -2161 1209 -2095
rect 1238 -2161 1242 -2095
rect 1262 -2161 1266 -2095
rect 1313 -2161 1317 -2095
rect 1205 -2172 1209 -2169
rect 1238 -2172 1242 -2169
rect 1262 -2172 1266 -2169
rect 1313 -2172 1317 -2169
rect 261 -2196 265 -2193
rect 677 -2196 681 -2193
rect 1121 -2196 1125 -2193
rect -575 -2224 -571 -2221
rect -554 -2224 -550 -2221
rect -509 -2224 -505 -2221
rect 357 -2224 361 -2221
rect 390 -2224 394 -2221
rect 414 -2224 418 -2221
rect 465 -2224 469 -2221
rect 1223 -2224 1227 -2221
rect 1256 -2224 1260 -2221
rect 1280 -2224 1284 -2221
rect 1331 -2224 1335 -2221
rect 59 -2228 63 -2225
rect -575 -2269 -571 -2232
rect -554 -2269 -550 -2232
rect -509 -2269 -505 -2232
rect 80 -2233 84 -2225
rect 125 -2228 129 -2225
rect 261 -2232 265 -2229
rect -30 -2257 -26 -2254
rect -575 -2280 -571 -2277
rect -554 -2280 -550 -2277
rect -509 -2280 -505 -2277
rect -30 -2296 -26 -2265
rect 261 -2277 265 -2240
rect 60 -2288 64 -2285
rect 81 -2288 85 -2285
rect 126 -2288 130 -2285
rect 261 -2288 265 -2285
rect -30 -2307 -26 -2304
rect -575 -2316 -571 -2313
rect -554 -2316 -550 -2313
rect -509 -2316 -505 -2313
rect -575 -2361 -571 -2324
rect -554 -2361 -550 -2324
rect -509 -2361 -505 -2324
rect 60 -2333 64 -2296
rect 81 -2333 85 -2296
rect 126 -2333 130 -2296
rect 357 -2298 361 -2232
rect 390 -2298 394 -2232
rect 414 -2298 418 -2232
rect 465 -2298 469 -2232
rect 1120 -2232 1124 -2229
rect 773 -2252 777 -2249
rect 806 -2252 810 -2249
rect 830 -2252 834 -2249
rect 881 -2252 885 -2249
rect 670 -2260 674 -2257
rect 670 -2305 674 -2268
rect 357 -2309 361 -2306
rect 390 -2309 394 -2306
rect 414 -2309 418 -2306
rect 465 -2309 469 -2306
rect 553 -2309 557 -2306
rect 574 -2309 578 -2306
rect 619 -2309 623 -2306
rect 670 -2316 674 -2313
rect 60 -2344 64 -2341
rect 81 -2349 85 -2341
rect 126 -2344 130 -2341
rect 553 -2354 557 -2317
rect 574 -2354 578 -2317
rect 619 -2354 623 -2317
rect 773 -2326 777 -2260
rect 806 -2326 810 -2260
rect 830 -2326 834 -2260
rect 881 -2326 885 -2260
rect 962 -2270 966 -2267
rect 983 -2270 987 -2267
rect 1028 -2270 1032 -2267
rect 1120 -2277 1124 -2240
rect 962 -2315 966 -2278
rect 983 -2315 987 -2278
rect 1028 -2315 1032 -2278
rect 1120 -2288 1124 -2285
rect 1223 -2298 1227 -2232
rect 1256 -2298 1260 -2232
rect 1280 -2298 1284 -2232
rect 1331 -2298 1335 -2232
rect 1443 -2265 1447 -2262
rect 1472 -2265 1476 -2262
rect 1496 -2265 1500 -2262
rect 1520 -2265 1524 -2262
rect 1567 -2265 1571 -2262
rect 1223 -2309 1227 -2306
rect 1256 -2309 1260 -2306
rect 1280 -2309 1284 -2306
rect 1331 -2309 1335 -2306
rect 962 -2326 966 -2323
rect 983 -2326 987 -2323
rect 1028 -2326 1032 -2323
rect 1443 -2327 1447 -2273
rect 1472 -2327 1476 -2273
rect 1496 -2327 1500 -2273
rect 1520 -2327 1524 -2273
rect 1567 -2327 1571 -2273
rect 773 -2337 777 -2334
rect 806 -2337 810 -2334
rect 830 -2337 834 -2334
rect 881 -2337 885 -2334
rect 1443 -2338 1447 -2335
rect 1472 -2338 1476 -2335
rect 1496 -2338 1500 -2335
rect 1520 -2338 1524 -2335
rect 1567 -2338 1571 -2335
rect 553 -2365 557 -2362
rect 574 -2365 578 -2362
rect 619 -2365 623 -2362
rect -575 -2372 -571 -2369
rect -554 -2372 -550 -2369
rect -509 -2372 -505 -2369
rect 41 -2466 45 -2463
rect 62 -2466 66 -2463
rect 83 -2466 87 -2463
rect 104 -2466 108 -2463
rect 172 -2466 176 -2463
rect 311 -2466 315 -2463
rect 332 -2466 336 -2463
rect 353 -2466 357 -2463
rect 374 -2466 378 -2463
rect 442 -2466 446 -2463
rect 41 -2534 45 -2474
rect 62 -2534 66 -2474
rect 83 -2534 87 -2474
rect 104 -2534 108 -2474
rect 172 -2534 176 -2474
rect 311 -2537 315 -2474
rect 332 -2537 336 -2474
rect 353 -2537 357 -2474
rect 374 -2537 378 -2474
rect 442 -2537 446 -2474
rect 41 -2545 45 -2542
rect 62 -2545 66 -2542
rect 83 -2545 87 -2542
rect 104 -2545 108 -2542
rect 172 -2545 176 -2542
rect 311 -2548 315 -2545
rect 332 -2548 336 -2545
rect 353 -2548 357 -2545
rect 374 -2548 378 -2545
rect 442 -2548 446 -2545
rect -574 -2600 -570 -2597
rect -553 -2600 -549 -2597
rect -508 -2600 -504 -2597
rect -574 -2645 -570 -2608
rect -553 -2645 -549 -2608
rect -508 -2645 -504 -2608
rect -574 -2656 -570 -2653
rect -553 -2656 -549 -2653
rect -508 -2656 -504 -2653
rect -577 -2692 -573 -2689
rect -556 -2692 -552 -2689
rect -511 -2692 -507 -2689
rect -577 -2737 -573 -2700
rect -556 -2737 -552 -2700
rect -511 -2737 -507 -2700
rect -577 -2748 -573 -2745
rect -556 -2748 -552 -2745
rect -511 -2748 -507 -2745
rect -76 -2759 -72 -2756
rect -55 -2759 -51 -2756
rect -10 -2759 -6 -2756
rect -577 -2784 -573 -2781
rect -556 -2784 -552 -2781
rect -511 -2784 -507 -2781
rect -577 -2829 -573 -2792
rect -556 -2829 -552 -2792
rect -511 -2829 -507 -2792
rect -76 -2804 -72 -2767
rect -55 -2804 -51 -2767
rect -10 -2804 -6 -2767
rect -76 -2815 -72 -2812
rect -55 -2815 -51 -2812
rect -10 -2815 -6 -2812
rect -577 -2840 -573 -2837
rect -556 -2840 -552 -2837
rect -511 -2840 -507 -2837
rect -76 -2852 -72 -2849
rect -55 -2852 -51 -2849
rect -10 -2852 -6 -2849
rect -577 -2876 -573 -2873
rect -556 -2876 -552 -2873
rect -511 -2876 -507 -2873
rect -577 -2921 -573 -2884
rect -556 -2921 -552 -2884
rect -511 -2921 -507 -2884
rect -76 -2897 -72 -2860
rect -55 -2897 -51 -2860
rect -10 -2897 -6 -2860
rect -76 -2908 -72 -2905
rect -55 -2908 -51 -2905
rect -10 -2908 -6 -2905
rect -577 -2932 -573 -2929
rect -556 -2932 -552 -2929
rect -511 -2932 -507 -2929
rect -76 -2944 -72 -2941
rect -55 -2944 -51 -2941
rect -10 -2944 -6 -2941
rect -572 -2967 -568 -2964
rect -551 -2967 -547 -2964
rect -506 -2967 -502 -2964
rect -572 -3012 -568 -2975
rect -551 -3012 -547 -2975
rect -506 -3012 -502 -2975
rect -76 -2989 -72 -2952
rect -55 -2989 -51 -2952
rect -10 -2989 -6 -2952
rect -76 -3000 -72 -2997
rect -55 -3000 -51 -2997
rect -10 -3000 -6 -2997
rect -572 -3023 -568 -3020
rect -551 -3023 -547 -3020
rect -506 -3023 -502 -3020
rect -76 -3037 -72 -3034
rect -55 -3037 -51 -3034
rect -10 -3037 -6 -3034
rect -575 -3059 -571 -3056
rect -554 -3059 -550 -3056
rect -509 -3059 -505 -3056
rect -575 -3104 -571 -3067
rect -554 -3104 -550 -3067
rect -509 -3104 -505 -3067
rect -76 -3082 -72 -3045
rect -55 -3082 -51 -3045
rect -10 -3082 -6 -3045
rect -76 -3093 -72 -3090
rect -55 -3093 -51 -3090
rect -10 -3093 -6 -3090
rect -575 -3115 -571 -3112
rect -554 -3115 -550 -3112
rect -509 -3115 -505 -3112
rect -575 -3151 -571 -3148
rect -554 -3151 -550 -3148
rect -509 -3151 -505 -3148
rect -575 -3196 -571 -3159
rect -554 -3196 -550 -3159
rect -509 -3196 -505 -3159
rect -575 -3207 -571 -3204
rect -554 -3207 -550 -3204
rect -509 -3207 -505 -3204
rect -575 -3243 -571 -3240
rect -554 -3243 -550 -3240
rect -509 -3243 -505 -3240
rect -575 -3288 -571 -3251
rect -554 -3288 -550 -3251
rect -509 -3288 -505 -3251
rect -575 -3299 -571 -3296
rect -554 -3299 -550 -3296
rect -509 -3299 -505 -3296
<< polycontact >>
rect -876 120 -872 124
rect -800 120 -796 124
rect -779 108 -775 112
rect -734 116 -730 120
rect -630 120 -626 124
rect -609 108 -605 112
rect -564 116 -560 120
rect -873 11 -869 15
rect -800 11 -796 15
rect -779 -1 -775 3
rect -734 7 -730 11
rect -634 11 -630 15
rect -613 -1 -609 3
rect -568 7 -564 11
rect -440 11 -436 15
rect -151 -43 -147 -39
rect 447 -43 451 -39
rect 1326 -43 1330 -39
rect 2094 -43 2098 -39
rect -224 -91 -220 -87
rect -130 -77 -126 -73
rect 374 -91 378 -87
rect -50 -111 -46 -107
rect -203 -125 -199 -121
rect -578 -144 -574 -140
rect -557 -156 -553 -152
rect -512 -148 -508 -144
rect 468 -77 472 -73
rect 1253 -91 1257 -87
rect 548 -111 552 -107
rect 395 -125 399 -121
rect -136 -152 -132 -148
rect 1347 -77 1351 -73
rect 2021 -91 2025 -87
rect 1427 -111 1431 -107
rect 1274 -125 1278 -121
rect -29 -145 -25 -141
rect 462 -152 466 -148
rect 2115 -77 2119 -73
rect 2195 -111 2199 -107
rect 2042 -125 2046 -121
rect 569 -145 573 -141
rect 1341 -152 1345 -148
rect 1448 -145 1452 -141
rect 2109 -152 2113 -148
rect 2216 -145 2220 -141
rect -115 -186 -111 -182
rect 483 -186 487 -182
rect 1362 -186 1366 -182
rect 2130 -186 2134 -182
rect -581 -236 -577 -232
rect -560 -248 -556 -244
rect -515 -240 -511 -236
rect -581 -328 -577 -324
rect -560 -340 -556 -336
rect -515 -332 -511 -328
rect 130 -346 134 -342
rect 873 -349 877 -345
rect 1632 -349 1636 -345
rect 2368 -349 2372 -345
rect -180 -394 -176 -390
rect -581 -420 -577 -416
rect -560 -432 -556 -428
rect -515 -424 -511 -420
rect 57 -394 61 -390
rect 151 -380 155 -376
rect 231 -414 235 -410
rect -253 -439 -249 -435
rect -159 -428 -155 -424
rect 78 -428 82 -424
rect 563 -397 567 -393
rect 800 -397 804 -393
rect 894 -383 898 -379
rect 1322 -397 1326 -393
rect 974 -417 978 -413
rect -79 -462 -75 -458
rect -232 -476 -228 -472
rect 145 -455 149 -451
rect 252 -448 256 -444
rect 490 -445 494 -441
rect 584 -431 588 -427
rect 821 -431 825 -427
rect 1559 -397 1563 -393
rect 1653 -383 1657 -379
rect 2058 -397 2062 -393
rect 1733 -417 1737 -413
rect 664 -465 668 -461
rect -576 -511 -572 -507
rect -555 -523 -551 -519
rect -510 -515 -506 -511
rect -165 -503 -161 -499
rect 511 -479 515 -475
rect -58 -496 -54 -492
rect 166 -489 170 -485
rect 888 -458 892 -454
rect 995 -451 999 -447
rect 1249 -445 1253 -441
rect 1343 -431 1347 -427
rect 1580 -431 1584 -427
rect 2295 -397 2299 -393
rect 2389 -383 2393 -379
rect 2469 -417 2473 -413
rect 1423 -465 1427 -461
rect 578 -506 582 -502
rect 1270 -479 1274 -475
rect 685 -499 689 -495
rect 909 -492 913 -488
rect 1647 -458 1651 -454
rect 1754 -451 1758 -447
rect 1985 -445 1989 -441
rect 2079 -431 2083 -427
rect 2316 -431 2320 -427
rect 2159 -465 2163 -461
rect 1337 -506 1341 -502
rect 2006 -479 2010 -475
rect 1444 -499 1448 -495
rect 1668 -492 1672 -488
rect 2383 -458 2387 -454
rect 2490 -451 2494 -447
rect 2073 -506 2077 -502
rect 2180 -499 2184 -495
rect 2404 -492 2408 -488
rect -144 -537 -140 -533
rect 599 -540 603 -536
rect 117 -561 121 -557
rect 138 -573 142 -569
rect 183 -565 187 -561
rect 276 -562 280 -558
rect -579 -603 -575 -599
rect -558 -615 -554 -611
rect -513 -607 -509 -603
rect 297 -570 301 -566
rect 344 -578 348 -574
rect 1358 -540 1362 -536
rect 2094 -540 2098 -536
rect 860 -564 864 -560
rect 881 -576 885 -572
rect 926 -568 930 -564
rect 1019 -565 1023 -561
rect -194 -612 -190 -608
rect -173 -624 -169 -620
rect -128 -616 -124 -612
rect 1040 -573 1044 -569
rect 1087 -581 1091 -577
rect 1619 -564 1623 -560
rect 1640 -576 1644 -572
rect 1685 -568 1689 -564
rect 1778 -565 1782 -561
rect 1799 -573 1803 -569
rect 1846 -581 1850 -577
rect 2355 -564 2359 -560
rect 2376 -576 2380 -572
rect 2421 -568 2425 -564
rect 2514 -565 2518 -561
rect 2535 -573 2539 -569
rect 2582 -581 2586 -577
rect 549 -615 553 -611
rect 570 -627 574 -623
rect 615 -619 619 -615
rect 1308 -615 1312 -611
rect 1329 -627 1333 -623
rect 1374 -619 1378 -615
rect 2044 -615 2048 -611
rect 2065 -627 2069 -623
rect 2110 -619 2114 -615
rect -579 -695 -575 -691
rect -558 -707 -554 -703
rect -513 -699 -509 -695
rect -579 -787 -575 -783
rect -558 -799 -554 -795
rect -513 -791 -509 -787
rect -122 -836 -118 -832
rect 476 -836 480 -832
rect 1355 -836 1359 -832
rect 2123 -836 2127 -832
rect -195 -884 -191 -880
rect -101 -870 -97 -866
rect 403 -884 407 -880
rect -21 -904 -17 -900
rect -174 -918 -170 -914
rect -578 -937 -574 -933
rect -557 -949 -553 -945
rect -512 -941 -508 -937
rect 497 -870 501 -866
rect 1282 -884 1286 -880
rect 577 -904 581 -900
rect 424 -918 428 -914
rect -107 -945 -103 -941
rect 1376 -870 1380 -866
rect 2050 -884 2054 -880
rect 1456 -904 1460 -900
rect 1303 -918 1307 -914
rect 0 -938 4 -934
rect 491 -945 495 -941
rect 2144 -870 2148 -866
rect 2224 -904 2228 -900
rect 2071 -918 2075 -914
rect 598 -938 602 -934
rect 1370 -945 1374 -941
rect 1477 -938 1481 -934
rect 2138 -945 2142 -941
rect 2245 -938 2249 -934
rect -86 -979 -82 -975
rect 512 -979 516 -975
rect 1391 -979 1395 -975
rect 2159 -979 2163 -975
rect -581 -1029 -577 -1025
rect -560 -1041 -556 -1037
rect -515 -1033 -511 -1029
rect -581 -1121 -577 -1117
rect -560 -1133 -556 -1129
rect -515 -1125 -511 -1121
rect 159 -1139 163 -1135
rect 902 -1142 906 -1138
rect 1661 -1142 1665 -1138
rect 2397 -1142 2401 -1138
rect -151 -1187 -147 -1183
rect -581 -1213 -577 -1209
rect -560 -1225 -556 -1221
rect -515 -1217 -511 -1213
rect 86 -1187 90 -1183
rect 180 -1173 184 -1169
rect 260 -1207 264 -1203
rect -224 -1232 -220 -1228
rect -130 -1221 -126 -1217
rect 107 -1221 111 -1217
rect 592 -1190 596 -1186
rect 829 -1190 833 -1186
rect 923 -1176 927 -1172
rect 1351 -1190 1355 -1186
rect 1003 -1210 1007 -1206
rect -50 -1255 -46 -1251
rect -203 -1269 -199 -1265
rect 174 -1248 178 -1244
rect 281 -1241 285 -1237
rect 519 -1238 523 -1234
rect 613 -1224 617 -1220
rect 850 -1224 854 -1220
rect 1588 -1190 1592 -1186
rect 1682 -1176 1686 -1172
rect 2087 -1190 2091 -1186
rect 1762 -1210 1766 -1206
rect 693 -1258 697 -1254
rect -576 -1304 -572 -1300
rect -555 -1316 -551 -1312
rect -510 -1308 -506 -1304
rect -136 -1296 -132 -1292
rect 540 -1272 544 -1268
rect -29 -1289 -25 -1285
rect 195 -1282 199 -1278
rect 917 -1251 921 -1247
rect 1024 -1244 1028 -1240
rect 1278 -1238 1282 -1234
rect 1372 -1224 1376 -1220
rect 1609 -1224 1613 -1220
rect 2324 -1190 2328 -1186
rect 2418 -1176 2422 -1172
rect 2498 -1210 2502 -1206
rect 1452 -1258 1456 -1254
rect 607 -1299 611 -1295
rect 1299 -1272 1303 -1268
rect 714 -1292 718 -1288
rect 938 -1285 942 -1281
rect 1676 -1251 1680 -1247
rect 1783 -1244 1787 -1240
rect 2014 -1238 2018 -1234
rect 2108 -1224 2112 -1220
rect 2345 -1224 2349 -1220
rect 2188 -1258 2192 -1254
rect 1366 -1299 1370 -1295
rect 2035 -1272 2039 -1268
rect 1473 -1292 1477 -1288
rect 1697 -1285 1701 -1281
rect 2412 -1251 2416 -1247
rect 2519 -1244 2523 -1240
rect 2102 -1299 2106 -1295
rect 2209 -1292 2213 -1288
rect 2433 -1285 2437 -1281
rect -115 -1330 -111 -1326
rect 628 -1333 632 -1329
rect 146 -1354 150 -1350
rect 167 -1366 171 -1362
rect 212 -1358 216 -1354
rect 305 -1355 309 -1351
rect -579 -1396 -575 -1392
rect -558 -1408 -554 -1404
rect -513 -1400 -509 -1396
rect 326 -1363 330 -1359
rect 373 -1371 377 -1367
rect 1387 -1333 1391 -1329
rect 2123 -1333 2127 -1329
rect 889 -1357 893 -1353
rect 910 -1369 914 -1365
rect 955 -1361 959 -1357
rect 1048 -1358 1052 -1354
rect -165 -1405 -161 -1401
rect -144 -1417 -140 -1413
rect -99 -1409 -95 -1405
rect 1069 -1366 1073 -1362
rect 1116 -1374 1120 -1370
rect 1648 -1357 1652 -1353
rect 1669 -1369 1673 -1365
rect 1714 -1361 1718 -1357
rect 1807 -1358 1811 -1354
rect 1828 -1366 1832 -1362
rect 1875 -1374 1879 -1370
rect 2384 -1357 2388 -1353
rect 2405 -1369 2409 -1365
rect 2450 -1361 2454 -1357
rect 2543 -1358 2547 -1354
rect 2564 -1366 2568 -1362
rect 2611 -1374 2615 -1370
rect 578 -1408 582 -1404
rect 599 -1420 603 -1416
rect 644 -1412 648 -1408
rect 1337 -1408 1341 -1404
rect 1358 -1420 1362 -1416
rect 1403 -1412 1407 -1408
rect 2073 -1408 2077 -1404
rect 2094 -1420 2098 -1416
rect 2139 -1412 2143 -1408
rect -579 -1488 -575 -1484
rect -558 -1500 -554 -1496
rect -513 -1492 -509 -1488
rect -579 -1580 -575 -1576
rect -558 -1592 -554 -1588
rect -513 -1584 -509 -1580
rect -578 -1700 -574 -1696
rect -557 -1712 -553 -1708
rect -512 -1704 -508 -1700
rect 15 -1756 19 -1752
rect -581 -1792 -577 -1788
rect -560 -1804 -556 -1800
rect -515 -1796 -511 -1792
rect 504 -1756 508 -1752
rect 888 -1756 892 -1752
rect -58 -1804 -54 -1800
rect 36 -1790 40 -1786
rect 116 -1824 120 -1820
rect -37 -1838 -33 -1834
rect 431 -1808 435 -1800
rect 242 -1828 246 -1824
rect 525 -1790 529 -1786
rect 1303 -1780 1307 -1776
rect 605 -1824 609 -1820
rect 452 -1838 456 -1834
rect 30 -1865 34 -1861
rect -581 -1884 -577 -1880
rect -560 -1896 -556 -1892
rect -515 -1888 -511 -1884
rect 815 -1808 819 -1800
rect 678 -1828 682 -1824
rect 909 -1790 913 -1786
rect 1023 -1824 1027 -1820
rect 836 -1838 840 -1834
rect 137 -1858 141 -1854
rect 519 -1865 523 -1861
rect 1096 -1828 1100 -1824
rect 1230 -1828 1234 -1824
rect 626 -1858 630 -1854
rect 903 -1865 907 -1861
rect 1324 -1814 1328 -1810
rect 1044 -1858 1048 -1854
rect 1404 -1848 1408 -1844
rect 1251 -1862 1255 -1858
rect 1472 -1852 1476 -1848
rect 1318 -1889 1322 -1885
rect 51 -1899 55 -1895
rect 540 -1899 544 -1895
rect 924 -1899 928 -1895
rect 1425 -1882 1429 -1878
rect 1339 -1923 1343 -1919
rect -581 -1976 -577 -1972
rect -560 -1988 -556 -1984
rect -515 -1980 -511 -1976
rect -576 -2067 -572 -2063
rect -555 -2079 -551 -2075
rect -510 -2071 -506 -2067
rect 335 -2111 339 -2107
rect -579 -2159 -575 -2155
rect -558 -2171 -554 -2167
rect -513 -2163 -509 -2159
rect 257 -2171 261 -2167
rect -32 -2191 -28 -2187
rect 55 -2199 59 -2195
rect 121 -2203 125 -2199
rect 368 -2119 372 -2115
rect 392 -2131 396 -2127
rect 443 -2147 447 -2143
rect 751 -2111 755 -2107
rect 673 -2171 677 -2167
rect 784 -2119 788 -2115
rect 808 -2131 812 -2127
rect 859 -2147 863 -2143
rect 1201 -2111 1205 -2107
rect 1117 -2171 1121 -2167
rect 1234 -2119 1238 -2115
rect 1258 -2131 1262 -2127
rect 1309 -2147 1313 -2143
rect -579 -2251 -575 -2247
rect -558 -2263 -554 -2259
rect -513 -2255 -509 -2251
rect 76 -2233 80 -2229
rect -34 -2288 -30 -2284
rect 257 -2266 261 -2262
rect 353 -2248 357 -2244
rect 56 -2315 60 -2311
rect -579 -2343 -575 -2339
rect -558 -2355 -554 -2351
rect -513 -2347 -509 -2343
rect 122 -2319 126 -2315
rect 386 -2256 390 -2252
rect 410 -2268 414 -2264
rect 461 -2284 465 -2280
rect 666 -2294 670 -2290
rect 769 -2276 773 -2272
rect 549 -2336 553 -2332
rect 77 -2349 81 -2345
rect 570 -2348 574 -2344
rect 615 -2340 619 -2336
rect 802 -2284 806 -2280
rect 826 -2296 830 -2292
rect 877 -2312 881 -2308
rect 1116 -2263 1120 -2259
rect 1219 -2248 1223 -2244
rect 958 -2297 962 -2293
rect 979 -2309 983 -2305
rect 1024 -2301 1028 -2297
rect 1252 -2256 1256 -2252
rect 1276 -2268 1280 -2264
rect 1327 -2284 1331 -2280
rect 1439 -2289 1443 -2285
rect 1468 -2305 1472 -2301
rect 1492 -2314 1496 -2310
rect 1516 -2323 1520 -2319
rect 1563 -2297 1567 -2293
rect 37 -2490 41 -2486
rect 58 -2498 62 -2494
rect 79 -2506 83 -2502
rect 100 -2514 104 -2510
rect 168 -2522 172 -2518
rect 307 -2490 311 -2486
rect 328 -2499 332 -2495
rect 349 -2508 353 -2504
rect 370 -2517 374 -2513
rect 438 -2525 442 -2521
rect -578 -2627 -574 -2623
rect -557 -2639 -553 -2635
rect -512 -2631 -508 -2627
rect -581 -2719 -577 -2715
rect -560 -2731 -556 -2727
rect -515 -2723 -511 -2719
rect -80 -2786 -76 -2782
rect -581 -2811 -577 -2807
rect -560 -2823 -556 -2819
rect -515 -2815 -511 -2811
rect -59 -2798 -55 -2794
rect -14 -2790 -10 -2786
rect -80 -2879 -76 -2875
rect -581 -2903 -577 -2899
rect -560 -2915 -556 -2911
rect -515 -2907 -511 -2903
rect -59 -2891 -55 -2887
rect -14 -2883 -10 -2879
rect -80 -2971 -76 -2967
rect -576 -2994 -572 -2990
rect -555 -3006 -551 -3002
rect -510 -2998 -506 -2994
rect -59 -2983 -55 -2979
rect -14 -2975 -10 -2971
rect -80 -3064 -76 -3060
rect -579 -3086 -575 -3082
rect -558 -3098 -554 -3094
rect -513 -3090 -509 -3086
rect -59 -3076 -55 -3072
rect -14 -3068 -10 -3064
rect -579 -3178 -575 -3174
rect -558 -3190 -554 -3186
rect -513 -3182 -509 -3178
rect -579 -3270 -575 -3266
rect -558 -3282 -554 -3278
rect -513 -3274 -509 -3270
<< metal1 >>
rect -920 188 -649 192
rect -920 86 -916 188
rect -906 180 -668 184
rect -906 124 -902 180
rect -891 163 -722 167
rect -877 145 -873 163
rect -801 145 -797 163
rect -768 145 -764 163
rect -735 145 -731 163
rect -906 120 -876 124
rect -867 120 -863 141
rect -804 120 -800 124
rect -791 120 -787 141
rect -867 116 -849 120
rect -791 116 -734 120
rect -867 106 -863 116
rect -877 86 -873 102
rect -920 82 -873 86
rect -853 86 -849 116
rect -820 108 -779 112
rect -820 86 -816 108
rect -768 100 -764 116
rect -725 115 -721 141
rect -725 111 -691 115
rect -725 100 -721 111
rect -853 82 -816 86
rect -801 86 -797 96
rect -735 86 -731 96
rect -801 82 -731 86
rect -904 -23 -900 82
rect -820 67 -816 82
rect -874 54 -722 58
rect -874 36 -870 54
rect -801 36 -797 54
rect -768 36 -764 54
rect -735 36 -731 54
rect -888 11 -873 15
rect -864 11 -860 32
rect -824 11 -800 15
rect -791 11 -787 32
rect -864 7 -846 11
rect -864 -3 -860 7
rect -791 7 -734 11
rect -815 -1 -779 3
rect -874 -23 -870 -7
rect -768 -9 -764 7
rect -725 6 -721 32
rect -725 2 -706 6
rect -725 -9 -721 2
rect -801 -23 -797 -13
rect -735 -23 -731 -13
rect -904 -27 -731 -23
rect -710 -81 -706 2
rect -941 -2570 -937 -89
rect -919 -85 -706 -81
rect -695 -81 -691 111
rect -672 112 -668 180
rect -653 159 -649 188
rect -638 163 -302 167
rect -631 145 -627 163
rect -598 145 -594 163
rect -565 145 -561 163
rect -634 120 -630 124
rect -621 120 -617 141
rect -621 116 -564 120
rect -672 108 -609 112
rect -672 3 -668 108
rect -598 100 -594 116
rect -555 115 -551 141
rect -555 111 -533 115
rect -555 100 -551 111
rect -631 86 -627 96
rect -565 86 -561 96
rect -638 82 -561 86
rect -659 54 -437 58
rect -635 36 -631 54
rect -602 36 -598 54
rect -569 36 -565 54
rect -441 36 -437 54
rect -638 11 -634 15
rect -625 11 -621 32
rect -625 7 -568 11
rect -672 -1 -613 3
rect -602 -9 -598 7
rect -559 6 -555 32
rect -431 15 -427 32
rect -444 11 -440 15
rect -431 11 -423 15
rect -306 12 -302 163
rect -559 2 -548 6
rect -559 -9 -555 2
rect -431 -10 -427 11
rect -635 -23 -631 -13
rect -569 -23 -565 -13
rect -306 8 -175 12
rect -441 -23 -437 -14
rect -638 -27 -437 -23
rect -569 -81 -565 -27
rect -695 -85 -604 -81
rect -569 -85 -325 -81
rect -919 -1643 -915 -85
rect -888 -3270 -884 -111
rect -868 -3178 -864 -111
rect -848 -3086 -844 -111
rect -828 -2994 -824 -111
rect -808 -2903 -804 -111
rect -788 -2811 -784 -111
rect -768 -2719 -764 -111
rect -748 -2627 -744 -111
rect -608 -152 -604 -85
rect -588 -101 -509 -97
rect -579 -119 -575 -101
rect -546 -119 -542 -101
rect -513 -119 -509 -101
rect -588 -144 -578 -140
rect -569 -144 -565 -123
rect -569 -148 -512 -144
rect -608 -156 -557 -152
rect -608 -244 -604 -156
rect -546 -164 -542 -148
rect -503 -149 -499 -123
rect -329 -124 -325 -85
rect -306 -142 -302 8
rect -179 4 -175 8
rect 399 9 414 13
rect 399 4 403 9
rect -183 0 403 4
rect 410 5 414 9
rect 1278 9 1293 13
rect 1278 4 1282 9
rect 415 0 1282 4
rect 1289 5 1293 9
rect 2046 8 2061 12
rect 2046 4 2050 8
rect 1294 0 2050 4
rect 2057 5 2061 8
rect 2062 0 2231 4
rect -244 -16 -171 -12
rect -244 -87 -240 -16
rect -175 -39 -171 -16
rect -152 -18 -148 0
rect -119 -18 -115 0
rect -175 -43 -151 -39
rect -142 -43 -138 -22
rect -142 -47 -74 -43
rect -225 -51 -188 -47
rect -225 -66 -221 -51
rect -192 -66 -188 -51
rect -119 -63 -115 -47
rect -248 -91 -224 -87
rect -215 -91 -211 -70
rect -134 -91 -130 -73
rect -215 -95 -130 -91
rect -192 -111 -188 -95
rect -503 -153 -478 -149
rect -503 -164 -499 -153
rect -579 -178 -575 -168
rect -513 -178 -509 -168
rect -207 -177 -203 -121
rect -162 -148 -158 -95
rect -144 -109 -96 -105
rect -78 -107 -74 -47
rect -51 -86 -47 0
rect -18 -86 -14 0
rect 354 -16 427 -12
rect -137 -127 -133 -109
rect -104 -127 -100 -109
rect -78 -111 -50 -107
rect -41 -111 -37 -90
rect 354 -87 358 -16
rect 423 -39 427 -16
rect 446 -18 450 0
rect 479 -18 483 0
rect 423 -43 447 -39
rect 456 -43 460 -22
rect 456 -47 524 -43
rect 373 -51 410 -47
rect 373 -66 377 -51
rect 406 -66 410 -51
rect 479 -63 483 -47
rect 350 -91 374 -87
rect 383 -91 387 -70
rect 464 -91 468 -73
rect 383 -95 468 -91
rect 406 -111 410 -95
rect -41 -115 7 -111
rect -18 -131 -14 -115
rect -162 -152 -136 -148
rect -127 -152 -123 -131
rect -33 -152 -29 -141
rect 391 -148 395 -121
rect -127 -156 -29 -152
rect 343 -152 395 -148
rect 436 -148 440 -95
rect 454 -109 502 -105
rect 520 -107 524 -47
rect 547 -86 551 0
rect 580 -1 1282 0
rect 580 -86 584 -1
rect 1233 -16 1306 -12
rect 461 -127 465 -109
rect 494 -127 498 -109
rect 520 -111 548 -107
rect 557 -111 561 -90
rect 1233 -87 1237 -16
rect 1302 -39 1306 -16
rect 1325 -18 1329 0
rect 1358 -18 1362 0
rect 1302 -43 1326 -39
rect 1335 -43 1339 -22
rect 1335 -47 1403 -43
rect 1252 -51 1289 -47
rect 1252 -66 1256 -51
rect 1285 -66 1289 -51
rect 1358 -63 1362 -47
rect 1229 -91 1253 -87
rect 1262 -91 1266 -70
rect 1343 -91 1347 -73
rect 1262 -95 1347 -91
rect 1285 -111 1289 -95
rect 557 -115 750 -111
rect 580 -131 584 -115
rect 436 -152 462 -148
rect 471 -152 475 -131
rect 565 -152 569 -141
rect 1270 -148 1274 -121
rect -104 -172 -100 -156
rect -579 -182 -509 -178
rect -392 -181 -203 -177
rect -588 -192 -512 -188
rect -582 -211 -578 -192
rect -549 -211 -545 -192
rect -516 -211 -512 -192
rect -588 -236 -581 -232
rect -572 -236 -568 -215
rect -572 -240 -515 -236
rect -608 -248 -560 -244
rect -608 -336 -604 -248
rect -549 -256 -545 -240
rect -506 -241 -502 -215
rect -412 -213 -400 -209
rect -506 -245 -469 -241
rect -506 -256 -502 -245
rect -582 -270 -578 -260
rect -516 -270 -512 -260
rect -582 -274 -512 -270
rect -588 -284 -512 -280
rect -582 -303 -578 -284
rect -549 -303 -545 -284
rect -516 -303 -512 -284
rect -588 -328 -581 -324
rect -572 -328 -568 -307
rect -572 -332 -515 -328
rect -608 -340 -560 -336
rect -608 -428 -604 -340
rect -549 -348 -545 -332
rect -506 -333 -502 -307
rect -506 -337 -461 -333
rect -506 -348 -502 -337
rect -582 -362 -578 -352
rect -516 -362 -512 -352
rect -582 -366 -512 -362
rect -588 -376 -512 -372
rect -582 -395 -578 -376
rect -549 -395 -545 -376
rect -516 -395 -512 -376
rect -588 -420 -581 -416
rect -572 -420 -568 -399
rect -572 -424 -515 -420
rect -608 -432 -560 -428
rect -608 -519 -604 -432
rect -549 -440 -545 -424
rect -506 -425 -502 -399
rect -506 -429 -494 -425
rect -506 -440 -502 -429
rect -498 -435 -494 -429
rect -498 -439 -453 -435
rect -582 -454 -578 -444
rect -516 -454 -512 -444
rect -582 -458 -512 -454
rect -586 -468 -507 -464
rect -577 -486 -573 -468
rect -544 -486 -540 -468
rect -511 -486 -507 -468
rect -586 -511 -576 -507
rect -567 -511 -563 -490
rect -567 -515 -510 -511
rect -608 -523 -555 -519
rect -608 -611 -604 -523
rect -544 -531 -540 -515
rect -501 -516 -497 -490
rect -444 -516 -440 -245
rect -501 -520 -440 -516
rect -501 -531 -497 -520
rect -577 -545 -573 -535
rect -511 -545 -507 -535
rect -577 -549 -507 -545
rect -586 -559 -510 -555
rect -580 -578 -576 -559
rect -547 -578 -543 -559
rect -514 -578 -510 -559
rect -586 -603 -579 -599
rect -570 -603 -566 -582
rect -570 -607 -513 -603
rect -608 -615 -558 -611
rect -608 -703 -604 -615
rect -547 -623 -543 -607
rect -504 -608 -500 -582
rect -430 -608 -426 -228
rect -504 -612 -426 -608
rect -504 -623 -500 -612
rect -580 -637 -576 -627
rect -514 -637 -510 -627
rect -580 -641 -510 -637
rect -586 -651 -510 -647
rect -580 -670 -576 -651
rect -547 -670 -543 -651
rect -514 -670 -510 -651
rect -586 -695 -579 -691
rect -570 -695 -566 -674
rect -570 -699 -513 -695
rect -608 -707 -558 -703
rect -608 -795 -604 -707
rect -547 -715 -543 -699
rect -504 -703 -500 -674
rect -412 -703 -408 -213
rect -504 -707 -408 -703
rect -504 -715 -500 -707
rect -580 -729 -576 -719
rect -514 -729 -510 -719
rect -580 -733 -510 -729
rect -586 -743 -510 -739
rect -580 -762 -576 -743
rect -547 -762 -543 -743
rect -514 -762 -510 -743
rect -586 -787 -579 -783
rect -570 -787 -566 -766
rect -570 -791 -513 -787
rect -608 -799 -558 -795
rect -547 -807 -543 -791
rect -504 -792 -500 -766
rect -392 -792 -388 -181
rect -207 -201 -203 -181
rect -119 -201 -115 -182
rect -207 -205 -115 -201
rect 343 -209 347 -152
rect 471 -156 569 -152
rect 1223 -156 1274 -148
rect 1315 -148 1319 -95
rect 1333 -109 1381 -105
rect 1399 -107 1403 -47
rect 1426 -86 1430 0
rect 1459 -86 1463 0
rect 1988 -1 1997 0
rect 2001 -16 2074 -12
rect 1340 -127 1344 -109
rect 1373 -127 1377 -109
rect 1399 -111 1427 -107
rect 1436 -111 1440 -90
rect 2001 -87 2005 -16
rect 2070 -39 2074 -16
rect 2093 -18 2097 0
rect 2126 -18 2130 0
rect 2070 -43 2094 -39
rect 2103 -43 2107 -22
rect 2103 -47 2171 -43
rect 2020 -51 2057 -47
rect 2020 -66 2024 -51
rect 2053 -66 2057 -51
rect 2126 -63 2130 -47
rect 1997 -91 2021 -87
rect 2030 -91 2034 -70
rect 2111 -91 2115 -73
rect 2030 -95 2115 -91
rect 2053 -111 2057 -95
rect 1436 -115 1520 -111
rect 1459 -131 1463 -115
rect 1315 -152 1341 -148
rect 1350 -152 1354 -131
rect 1444 -152 1448 -141
rect 2038 -148 2042 -121
rect 1350 -156 1448 -152
rect 1984 -156 2042 -148
rect 2083 -148 2087 -95
rect 2101 -109 2149 -105
rect 2167 -107 2171 -47
rect 2194 -86 2198 0
rect 2227 -86 2231 0
rect 2108 -127 2112 -109
rect 2141 -127 2145 -109
rect 2167 -111 2195 -107
rect 2204 -111 2208 -90
rect 2204 -115 2254 -111
rect 2227 -131 2231 -115
rect 2083 -152 2109 -148
rect 2118 -152 2122 -131
rect 2212 -152 2216 -141
rect 2118 -156 2216 -152
rect 494 -172 498 -156
rect 479 -209 483 -182
rect -238 -213 483 -209
rect 1223 -228 1227 -156
rect 1270 -201 1274 -156
rect 1373 -172 1377 -156
rect 1358 -201 1362 -182
rect 1270 -205 1362 -201
rect -238 -232 1227 -228
rect 1984 -245 1988 -156
rect 2038 -201 2042 -156
rect 2141 -172 2145 -156
rect 2126 -201 2130 -182
rect 2038 -205 2130 -201
rect -238 -249 1988 -245
rect 98 -303 298 -299
rect 33 -319 110 -315
rect -212 -351 -12 -347
rect -277 -367 -200 -363
rect -277 -434 -273 -367
rect -204 -390 -200 -367
rect -181 -369 -177 -351
rect -148 -369 -144 -351
rect -204 -394 -180 -390
rect -171 -394 -167 -373
rect -171 -398 -103 -394
rect -254 -402 -217 -398
rect -254 -417 -250 -402
rect -221 -417 -217 -402
rect -148 -414 -144 -398
rect -272 -439 -253 -435
rect -277 -608 -273 -439
rect -244 -442 -240 -421
rect -163 -442 -159 -424
rect -244 -446 -159 -442
rect -221 -462 -217 -446
rect -236 -499 -232 -472
rect -252 -503 -232 -499
rect -191 -499 -187 -446
rect -173 -460 -125 -456
rect -107 -458 -103 -398
rect -80 -437 -76 -351
rect -47 -437 -43 -351
rect -166 -478 -162 -460
rect -133 -478 -129 -460
rect -107 -462 -79 -458
rect -70 -464 -66 -441
rect -70 -468 -27 -464
rect -47 -482 -43 -468
rect -191 -503 -165 -499
rect -156 -503 -152 -482
rect -62 -503 -58 -492
rect -236 -552 -232 -503
rect -156 -507 -58 -503
rect -133 -523 -129 -507
rect -148 -552 -144 -533
rect -236 -558 -144 -552
rect -16 -565 -12 -351
rect 33 -390 37 -319
rect 106 -342 110 -319
rect 129 -321 133 -303
rect 162 -321 166 -303
rect 106 -346 130 -342
rect 139 -346 143 -325
rect 139 -350 207 -346
rect 56 -354 93 -350
rect 56 -369 60 -354
rect 89 -369 93 -354
rect 162 -366 166 -350
rect 8 -394 57 -390
rect 66 -394 70 -373
rect 147 -394 151 -376
rect 33 -557 37 -394
rect 66 -398 151 -394
rect 89 -414 93 -398
rect 74 -451 78 -424
rect 58 -455 78 -451
rect 119 -451 123 -398
rect 137 -412 185 -408
rect 203 -410 207 -350
rect 230 -389 234 -303
rect 263 -389 267 -303
rect 294 -350 298 -303
rect 841 -306 1041 -302
rect 1600 -306 1800 -302
rect 2336 -306 2536 -302
rect 776 -322 853 -318
rect 294 -354 526 -350
rect 531 -354 731 -350
rect 144 -430 148 -412
rect 177 -430 181 -412
rect 203 -414 231 -410
rect 240 -414 244 -393
rect 240 -418 283 -414
rect 263 -434 267 -418
rect 119 -455 145 -451
rect 154 -455 158 -434
rect 248 -455 252 -444
rect 74 -504 78 -455
rect 154 -459 252 -455
rect 177 -475 181 -459
rect 162 -504 166 -485
rect 74 -508 166 -504
rect 294 -514 298 -354
rect 466 -370 543 -366
rect 466 -441 470 -370
rect 539 -393 543 -370
rect 562 -372 566 -354
rect 595 -372 599 -354
rect 539 -397 563 -393
rect 572 -397 576 -376
rect 572 -401 640 -397
rect 489 -405 526 -401
rect 489 -420 493 -405
rect 522 -420 526 -405
rect 595 -417 599 -401
rect 423 -445 490 -441
rect 499 -445 503 -424
rect 580 -445 584 -427
rect 116 -518 347 -514
rect 116 -536 120 -518
rect 149 -536 153 -518
rect 182 -536 186 -518
rect 275 -536 279 -518
rect 343 -536 347 -518
rect 33 -561 117 -557
rect 126 -561 130 -540
rect 192 -558 196 -540
rect 126 -565 183 -561
rect 192 -562 276 -558
rect -195 -569 -12 -565
rect -195 -587 -191 -569
rect -162 -587 -158 -569
rect -129 -587 -125 -569
rect 99 -573 138 -569
rect 149 -581 153 -565
rect 192 -581 196 -562
rect 272 -570 297 -566
rect 310 -574 314 -540
rect 353 -561 357 -540
rect 423 -561 427 -445
rect 353 -565 427 -561
rect 285 -578 344 -574
rect 285 -584 289 -578
rect 353 -584 357 -565
rect -277 -612 -194 -608
rect -185 -612 -181 -591
rect -185 -616 -128 -612
rect -211 -624 -173 -620
rect -162 -632 -158 -616
rect -119 -617 -115 -591
rect 116 -600 120 -585
rect 182 -600 186 -585
rect 275 -600 279 -588
rect 308 -600 312 -588
rect 343 -600 347 -588
rect 109 -604 347 -600
rect -119 -621 208 -617
rect -119 -632 -115 -621
rect -195 -648 -191 -636
rect -129 -648 -125 -636
rect -195 -652 -125 -648
rect 343 -651 347 -604
rect 466 -611 470 -445
rect 499 -449 584 -445
rect 522 -465 526 -449
rect 507 -502 511 -475
rect 491 -506 511 -502
rect 552 -502 556 -449
rect 570 -463 618 -459
rect 636 -461 640 -401
rect 663 -440 667 -354
rect 696 -440 700 -354
rect 577 -481 581 -463
rect 610 -481 614 -463
rect 636 -465 664 -461
rect 673 -467 677 -444
rect 673 -471 716 -467
rect 696 -485 700 -471
rect 552 -506 578 -502
rect 587 -506 591 -485
rect 681 -506 685 -495
rect 507 -555 511 -506
rect 587 -510 685 -506
rect 610 -526 614 -510
rect 595 -555 599 -536
rect 507 -559 599 -555
rect 727 -568 731 -354
rect 776 -393 780 -322
rect 849 -345 853 -322
rect 872 -324 876 -306
rect 905 -324 909 -306
rect 849 -349 873 -345
rect 882 -349 886 -328
rect 882 -353 950 -349
rect 799 -357 836 -353
rect 799 -372 803 -357
rect 832 -372 836 -357
rect 905 -369 909 -353
rect 751 -397 800 -393
rect 809 -397 813 -376
rect 890 -397 894 -379
rect 776 -560 780 -397
rect 809 -401 894 -397
rect 832 -417 836 -401
rect 817 -454 821 -427
rect 801 -458 821 -454
rect 862 -454 866 -401
rect 880 -415 928 -411
rect 946 -413 950 -353
rect 973 -392 977 -306
rect 1006 -392 1010 -306
rect 1037 -350 1041 -306
rect 1535 -322 1612 -318
rect 1037 -354 1285 -350
rect 1290 -354 1490 -350
rect 887 -433 891 -415
rect 920 -433 924 -415
rect 946 -417 974 -413
rect 983 -417 987 -396
rect 983 -421 1026 -417
rect 1006 -437 1010 -421
rect 862 -458 888 -454
rect 897 -458 901 -437
rect 991 -458 995 -447
rect 817 -507 821 -458
rect 897 -462 995 -458
rect 920 -478 924 -462
rect 905 -507 909 -488
rect 817 -511 909 -507
rect 1037 -517 1041 -354
rect 1225 -370 1302 -366
rect 1225 -441 1229 -370
rect 1298 -393 1302 -370
rect 1321 -372 1325 -354
rect 1354 -372 1358 -354
rect 1298 -397 1322 -393
rect 1331 -397 1335 -376
rect 1331 -401 1399 -397
rect 1248 -405 1285 -401
rect 1248 -420 1252 -405
rect 1281 -420 1285 -405
rect 1354 -417 1358 -401
rect 1176 -445 1249 -441
rect 1258 -445 1262 -424
rect 1339 -445 1343 -427
rect 859 -521 1090 -517
rect 859 -539 863 -521
rect 892 -539 896 -521
rect 925 -539 929 -521
rect 1018 -539 1022 -521
rect 1086 -539 1090 -521
rect 776 -564 860 -560
rect 869 -564 873 -543
rect 935 -561 939 -543
rect 869 -568 926 -564
rect 935 -565 1019 -561
rect 548 -572 731 -568
rect 548 -590 552 -572
rect 581 -590 585 -572
rect 614 -590 618 -572
rect 842 -576 881 -572
rect 892 -584 896 -568
rect 935 -584 939 -565
rect 1015 -573 1040 -569
rect 1053 -577 1057 -543
rect 1096 -564 1100 -543
rect 1176 -564 1180 -445
rect 1096 -568 1180 -564
rect 1028 -581 1087 -577
rect 1028 -587 1032 -581
rect 1096 -587 1100 -568
rect 466 -615 549 -611
rect 558 -615 562 -594
rect 558 -619 615 -615
rect 532 -627 570 -623
rect 581 -635 585 -619
rect 624 -620 628 -594
rect 859 -603 863 -588
rect 925 -603 929 -588
rect 1018 -603 1022 -591
rect 1051 -603 1055 -591
rect 1086 -603 1090 -591
rect 852 -607 1090 -603
rect 624 -624 951 -620
rect 624 -635 628 -624
rect 548 -651 552 -639
rect 614 -651 618 -639
rect 1086 -650 1090 -607
rect 1225 -611 1229 -445
rect 1258 -449 1343 -445
rect 1281 -465 1285 -449
rect 1266 -502 1270 -475
rect 1250 -506 1270 -502
rect 1311 -502 1315 -449
rect 1329 -463 1377 -459
rect 1395 -461 1399 -401
rect 1422 -440 1426 -354
rect 1455 -440 1459 -354
rect 1336 -481 1340 -463
rect 1369 -481 1373 -463
rect 1395 -465 1423 -461
rect 1432 -467 1436 -444
rect 1432 -471 1475 -467
rect 1455 -485 1459 -471
rect 1311 -506 1337 -502
rect 1346 -506 1350 -485
rect 1440 -506 1444 -495
rect 1266 -555 1270 -506
rect 1346 -510 1444 -506
rect 1369 -526 1373 -510
rect 1354 -555 1358 -536
rect 1266 -559 1358 -555
rect 1270 -561 1358 -559
rect 1486 -568 1490 -354
rect 1535 -393 1539 -322
rect 1608 -345 1612 -322
rect 1631 -324 1635 -306
rect 1664 -324 1668 -306
rect 1608 -349 1632 -345
rect 1641 -349 1645 -328
rect 1641 -353 1709 -349
rect 1558 -357 1595 -353
rect 1558 -372 1562 -357
rect 1591 -372 1595 -357
rect 1664 -369 1668 -353
rect 1535 -397 1559 -393
rect 1568 -397 1572 -376
rect 1649 -397 1653 -379
rect 1535 -560 1539 -397
rect 1568 -401 1653 -397
rect 1591 -417 1595 -401
rect 1576 -454 1580 -427
rect 1560 -458 1580 -454
rect 1621 -454 1625 -401
rect 1639 -415 1687 -411
rect 1705 -413 1709 -353
rect 1732 -392 1736 -306
rect 1765 -392 1769 -306
rect 1796 -350 1800 -306
rect 2271 -322 2348 -318
rect 1796 -354 2021 -350
rect 2026 -354 2226 -350
rect 1646 -433 1650 -415
rect 1679 -433 1683 -415
rect 1705 -417 1733 -413
rect 1742 -417 1746 -396
rect 1742 -421 1785 -417
rect 1765 -437 1769 -421
rect 1621 -458 1647 -454
rect 1656 -458 1660 -437
rect 1750 -458 1754 -447
rect 1576 -507 1580 -458
rect 1656 -462 1754 -458
rect 1679 -478 1683 -462
rect 1796 -484 1800 -354
rect 1961 -370 2038 -366
rect 1961 -441 1965 -370
rect 2034 -393 2038 -370
rect 2057 -372 2061 -354
rect 2090 -372 2094 -354
rect 2034 -397 2058 -393
rect 2067 -397 2071 -376
rect 2067 -401 2135 -397
rect 1984 -405 2021 -401
rect 1984 -420 1988 -405
rect 2017 -420 2021 -405
rect 2090 -417 2094 -401
rect 1770 -488 1800 -484
rect 1906 -445 1985 -441
rect 1994 -445 1998 -424
rect 2075 -445 2079 -427
rect 1664 -507 1668 -488
rect 1576 -511 1668 -507
rect 1770 -517 1774 -488
rect 1618 -521 1849 -517
rect 1618 -539 1622 -521
rect 1651 -539 1655 -521
rect 1684 -539 1688 -521
rect 1777 -539 1781 -521
rect 1845 -539 1849 -521
rect 1535 -564 1619 -560
rect 1628 -564 1632 -543
rect 1694 -561 1698 -543
rect 1628 -568 1685 -564
rect 1694 -565 1778 -561
rect 1307 -572 1490 -568
rect 1307 -590 1311 -572
rect 1340 -590 1344 -572
rect 1373 -590 1377 -572
rect 1601 -576 1640 -572
rect 1651 -584 1655 -568
rect 1694 -584 1698 -565
rect 1774 -573 1799 -569
rect 1812 -577 1816 -543
rect 1855 -564 1859 -543
rect 1906 -564 1910 -445
rect 1855 -568 1910 -564
rect 1787 -581 1846 -577
rect 1787 -587 1791 -581
rect 1855 -587 1859 -568
rect 1225 -615 1308 -611
rect 1317 -615 1321 -594
rect 1317 -619 1374 -615
rect 1291 -627 1329 -623
rect 1340 -635 1344 -619
rect 1383 -620 1387 -594
rect 1618 -603 1622 -588
rect 1684 -603 1688 -588
rect 1777 -603 1781 -591
rect 1810 -603 1814 -591
rect 1845 -603 1849 -591
rect 1611 -607 1849 -603
rect 1383 -624 1710 -620
rect 1383 -635 1387 -624
rect 1307 -650 1311 -639
rect 1373 -649 1377 -639
rect 343 -655 618 -651
rect 1086 -654 1372 -650
rect 1845 -650 1849 -607
rect 1961 -611 1965 -445
rect 1994 -449 2079 -445
rect 2017 -465 2021 -449
rect 2002 -502 2006 -475
rect 1986 -506 2006 -502
rect 2047 -502 2051 -449
rect 2065 -463 2113 -459
rect 2131 -461 2135 -401
rect 2158 -440 2162 -354
rect 2191 -440 2195 -354
rect 2072 -481 2076 -463
rect 2105 -481 2109 -463
rect 2131 -465 2159 -461
rect 2168 -467 2172 -444
rect 2168 -471 2211 -467
rect 2191 -485 2195 -471
rect 2047 -506 2073 -502
rect 2082 -506 2086 -485
rect 2176 -506 2180 -495
rect 2002 -555 2006 -506
rect 2082 -510 2180 -506
rect 2105 -526 2109 -510
rect 2090 -555 2094 -536
rect 2002 -559 2094 -555
rect 2006 -561 2094 -559
rect 2222 -568 2226 -354
rect 2271 -393 2275 -322
rect 2344 -345 2348 -322
rect 2367 -324 2371 -306
rect 2400 -324 2404 -306
rect 2344 -349 2368 -345
rect 2377 -349 2381 -328
rect 2377 -353 2445 -349
rect 2294 -357 2331 -353
rect 2294 -372 2298 -357
rect 2327 -372 2331 -357
rect 2400 -369 2404 -353
rect 2271 -397 2295 -393
rect 2304 -397 2308 -376
rect 2385 -397 2389 -379
rect 2271 -560 2275 -397
rect 2304 -401 2389 -397
rect 2327 -417 2331 -401
rect 2312 -454 2316 -427
rect 2296 -458 2316 -454
rect 2357 -454 2361 -401
rect 2375 -415 2423 -411
rect 2441 -413 2445 -353
rect 2468 -392 2472 -306
rect 2501 -392 2505 -306
rect 2382 -433 2386 -415
rect 2415 -433 2419 -415
rect 2441 -417 2469 -413
rect 2478 -417 2482 -396
rect 2478 -421 2521 -417
rect 2501 -437 2505 -421
rect 2357 -458 2383 -454
rect 2392 -458 2396 -437
rect 2486 -458 2490 -447
rect 2312 -507 2316 -458
rect 2392 -462 2490 -458
rect 2415 -478 2419 -462
rect 2532 -484 2536 -306
rect 2506 -488 2536 -484
rect 2400 -507 2404 -488
rect 2312 -511 2404 -507
rect 2506 -517 2510 -488
rect 2354 -521 2585 -517
rect 2354 -539 2358 -521
rect 2387 -539 2391 -521
rect 2420 -539 2424 -521
rect 2513 -539 2517 -521
rect 2581 -539 2585 -521
rect 2271 -564 2355 -560
rect 2364 -564 2368 -543
rect 2430 -561 2434 -543
rect 2364 -568 2421 -564
rect 2430 -565 2514 -561
rect 2043 -572 2226 -568
rect 2043 -590 2047 -572
rect 2076 -590 2080 -572
rect 2109 -590 2113 -572
rect 2337 -576 2376 -572
rect 2387 -584 2391 -568
rect 2430 -584 2434 -565
rect 2510 -573 2535 -569
rect 2548 -577 2552 -543
rect 2591 -564 2595 -543
rect 2591 -568 2603 -564
rect 2523 -581 2582 -577
rect 2523 -587 2527 -581
rect 2591 -587 2595 -568
rect 1961 -615 2044 -611
rect 2053 -615 2057 -594
rect 2053 -619 2110 -615
rect 2027 -627 2065 -623
rect 2076 -635 2080 -619
rect 2119 -620 2123 -594
rect 2354 -603 2358 -588
rect 2420 -603 2424 -588
rect 2513 -603 2517 -591
rect 2546 -603 2550 -591
rect 2581 -603 2585 -591
rect 2347 -607 2585 -603
rect 2119 -624 2446 -620
rect 2119 -635 2123 -624
rect 2043 -650 2047 -639
rect 2109 -648 2113 -639
rect 1845 -653 2108 -650
rect -274 -670 438 -666
rect 1212 -683 1216 -679
rect -274 -687 1216 -683
rect 1936 -695 1940 -690
rect -274 -699 1940 -695
rect -504 -796 -388 -792
rect -277 -785 -146 -781
rect -504 -807 -500 -796
rect -354 -808 -337 -804
rect -580 -821 -576 -811
rect -514 -821 -510 -811
rect -580 -825 -510 -821
rect -354 -844 -350 -808
rect -608 -848 -350 -844
rect -608 -884 -604 -848
rect -625 -888 -604 -884
rect -608 -945 -604 -888
rect -277 -890 -273 -785
rect -150 -789 -146 -785
rect 428 -784 443 -780
rect 428 -789 432 -784
rect -154 -793 432 -789
rect 439 -788 443 -784
rect 1307 -784 1322 -780
rect 1307 -789 1311 -784
rect 444 -793 1311 -789
rect 1318 -788 1322 -784
rect 2075 -785 2090 -781
rect 2075 -789 2079 -785
rect 1323 -793 2079 -789
rect 2086 -788 2090 -785
rect 2091 -793 2260 -789
rect -215 -809 -142 -805
rect -215 -880 -211 -809
rect -146 -832 -142 -809
rect -123 -811 -119 -793
rect -90 -811 -86 -793
rect -146 -836 -122 -832
rect -113 -836 -109 -815
rect -113 -840 -45 -836
rect -196 -844 -159 -840
rect -196 -859 -192 -844
rect -163 -859 -159 -844
rect -90 -856 -86 -840
rect -219 -884 -195 -880
rect -186 -884 -182 -863
rect -105 -884 -101 -866
rect -186 -888 -101 -884
rect -588 -894 -273 -890
rect -579 -912 -575 -894
rect -546 -912 -542 -894
rect -513 -912 -509 -894
rect -588 -937 -578 -933
rect -569 -937 -565 -916
rect -569 -941 -512 -937
rect -608 -949 -557 -945
rect -608 -1037 -604 -949
rect -546 -957 -542 -941
rect -503 -942 -499 -916
rect -399 -922 -321 -918
rect -277 -935 -273 -894
rect -163 -904 -159 -888
rect -503 -946 -478 -942
rect -503 -957 -499 -946
rect -579 -971 -575 -961
rect -513 -971 -509 -961
rect -178 -970 -174 -914
rect -133 -941 -129 -888
rect -115 -902 -67 -898
rect -49 -900 -45 -840
rect -22 -879 -18 -793
rect 11 -879 15 -793
rect 383 -809 456 -805
rect -108 -920 -104 -902
rect -75 -920 -71 -902
rect -49 -904 -21 -900
rect -12 -904 -8 -883
rect 383 -880 387 -809
rect 452 -832 456 -809
rect 475 -811 479 -793
rect 508 -811 512 -793
rect 452 -836 476 -832
rect 485 -836 489 -815
rect 485 -840 553 -836
rect 402 -844 439 -840
rect 402 -859 406 -844
rect 435 -859 439 -844
rect 508 -856 512 -840
rect 379 -884 403 -880
rect 412 -884 416 -863
rect 493 -884 497 -866
rect 412 -888 497 -884
rect 435 -904 439 -888
rect -12 -908 36 -904
rect 11 -924 15 -908
rect -133 -945 -107 -941
rect -98 -945 -94 -924
rect -4 -945 0 -934
rect 420 -941 424 -914
rect -98 -949 0 -945
rect 372 -945 424 -941
rect 465 -941 469 -888
rect 483 -902 531 -898
rect 549 -900 553 -840
rect 576 -879 580 -793
rect 609 -794 1311 -793
rect 609 -879 613 -794
rect 1262 -809 1335 -805
rect 490 -920 494 -902
rect 523 -920 527 -902
rect 549 -904 577 -900
rect 586 -904 590 -883
rect 1262 -880 1266 -809
rect 1331 -832 1335 -809
rect 1354 -811 1358 -793
rect 1387 -811 1391 -793
rect 1331 -836 1355 -832
rect 1364 -836 1368 -815
rect 1364 -840 1432 -836
rect 1281 -844 1318 -840
rect 1281 -859 1285 -844
rect 1314 -859 1318 -844
rect 1387 -856 1391 -840
rect 1258 -884 1282 -880
rect 1291 -884 1295 -863
rect 1372 -884 1376 -866
rect 1291 -888 1376 -884
rect 1314 -904 1318 -888
rect 586 -908 779 -904
rect 609 -924 613 -908
rect 465 -945 491 -941
rect 500 -945 504 -924
rect 594 -945 598 -934
rect 1299 -941 1303 -914
rect -75 -965 -71 -949
rect -579 -975 -509 -971
rect -392 -974 -174 -970
rect -588 -985 -512 -981
rect -582 -1004 -578 -985
rect -549 -1004 -545 -985
rect -516 -1004 -512 -985
rect -588 -1029 -581 -1025
rect -572 -1029 -568 -1008
rect -572 -1033 -515 -1029
rect -608 -1041 -560 -1037
rect -608 -1129 -604 -1041
rect -549 -1049 -545 -1033
rect -506 -1034 -502 -1008
rect -412 -1006 -400 -1002
rect -506 -1038 -469 -1034
rect -506 -1049 -502 -1038
rect -582 -1063 -578 -1053
rect -516 -1063 -512 -1053
rect -582 -1067 -512 -1063
rect -588 -1077 -512 -1073
rect -582 -1096 -578 -1077
rect -549 -1096 -545 -1077
rect -516 -1096 -512 -1077
rect -588 -1121 -581 -1117
rect -572 -1121 -568 -1100
rect -572 -1125 -515 -1121
rect -608 -1133 -560 -1129
rect -608 -1221 -604 -1133
rect -549 -1141 -545 -1125
rect -506 -1126 -502 -1100
rect -506 -1130 -461 -1126
rect -506 -1141 -502 -1130
rect -582 -1155 -578 -1145
rect -516 -1155 -512 -1145
rect -582 -1159 -512 -1155
rect -588 -1169 -512 -1165
rect -582 -1188 -578 -1169
rect -549 -1188 -545 -1169
rect -516 -1188 -512 -1169
rect -588 -1213 -581 -1209
rect -572 -1213 -568 -1192
rect -572 -1217 -515 -1213
rect -608 -1225 -560 -1221
rect -608 -1312 -604 -1225
rect -549 -1233 -545 -1217
rect -506 -1218 -502 -1192
rect -506 -1222 -494 -1218
rect -506 -1233 -502 -1222
rect -498 -1228 -494 -1222
rect -498 -1232 -453 -1228
rect -582 -1247 -578 -1237
rect -516 -1247 -512 -1237
rect -582 -1251 -512 -1247
rect -586 -1261 -507 -1257
rect -577 -1279 -573 -1261
rect -544 -1279 -540 -1261
rect -511 -1279 -507 -1261
rect -586 -1304 -576 -1300
rect -567 -1304 -563 -1283
rect -567 -1308 -510 -1304
rect -608 -1316 -555 -1312
rect -608 -1404 -604 -1316
rect -544 -1324 -540 -1308
rect -501 -1309 -497 -1283
rect -444 -1309 -440 -1038
rect -501 -1313 -440 -1309
rect -501 -1324 -497 -1313
rect -577 -1338 -573 -1328
rect -511 -1338 -507 -1328
rect -577 -1342 -507 -1338
rect -586 -1352 -510 -1348
rect -580 -1371 -576 -1352
rect -547 -1371 -543 -1352
rect -514 -1371 -510 -1352
rect -586 -1396 -579 -1392
rect -570 -1396 -566 -1375
rect -570 -1400 -513 -1396
rect -608 -1408 -558 -1404
rect -608 -1496 -604 -1408
rect -547 -1416 -543 -1400
rect -504 -1401 -500 -1375
rect -430 -1401 -426 -1021
rect -504 -1405 -426 -1401
rect -504 -1416 -500 -1405
rect -580 -1430 -576 -1420
rect -514 -1430 -510 -1420
rect -580 -1434 -510 -1430
rect -586 -1444 -510 -1440
rect -580 -1463 -576 -1444
rect -547 -1463 -543 -1444
rect -514 -1463 -510 -1444
rect -586 -1488 -579 -1484
rect -570 -1488 -566 -1467
rect -570 -1492 -513 -1488
rect -608 -1500 -558 -1496
rect -608 -1588 -604 -1500
rect -547 -1508 -543 -1492
rect -504 -1496 -500 -1467
rect -412 -1496 -408 -1006
rect -504 -1500 -408 -1496
rect -504 -1508 -500 -1500
rect -580 -1522 -576 -1512
rect -514 -1522 -510 -1512
rect -580 -1526 -510 -1522
rect -586 -1536 -510 -1532
rect -580 -1555 -576 -1536
rect -547 -1555 -543 -1536
rect -514 -1555 -510 -1536
rect -586 -1580 -579 -1576
rect -570 -1580 -566 -1559
rect -570 -1584 -513 -1580
rect -608 -1592 -558 -1588
rect -547 -1600 -543 -1584
rect -504 -1585 -500 -1559
rect -392 -1585 -388 -974
rect -178 -994 -174 -974
rect -90 -994 -86 -975
rect -178 -998 -86 -994
rect 372 -1002 376 -945
rect 500 -949 598 -945
rect 1252 -949 1303 -941
rect 1344 -941 1348 -888
rect 1362 -902 1410 -898
rect 1428 -900 1432 -840
rect 1455 -879 1459 -793
rect 1488 -879 1492 -793
rect 2017 -794 2026 -793
rect 2030 -809 2103 -805
rect 1369 -920 1373 -902
rect 1402 -920 1406 -902
rect 1428 -904 1456 -900
rect 1465 -904 1469 -883
rect 2030 -880 2034 -809
rect 2099 -832 2103 -809
rect 2122 -811 2126 -793
rect 2155 -811 2159 -793
rect 2099 -836 2123 -832
rect 2132 -836 2136 -815
rect 2132 -840 2200 -836
rect 2049 -844 2086 -840
rect 2049 -859 2053 -844
rect 2082 -859 2086 -844
rect 2155 -856 2159 -840
rect 2026 -884 2050 -880
rect 2059 -884 2063 -863
rect 2140 -884 2144 -866
rect 2059 -888 2144 -884
rect 2082 -904 2086 -888
rect 1465 -908 1549 -904
rect 1488 -924 1492 -908
rect 1344 -945 1370 -941
rect 1379 -945 1383 -924
rect 1473 -945 1477 -934
rect 2067 -941 2071 -914
rect 1379 -949 1477 -945
rect 2013 -949 2071 -941
rect 2112 -941 2116 -888
rect 2130 -902 2178 -898
rect 2196 -900 2200 -840
rect 2223 -879 2227 -793
rect 2256 -879 2260 -793
rect 2137 -920 2141 -902
rect 2170 -920 2174 -902
rect 2196 -904 2224 -900
rect 2233 -904 2237 -883
rect 2233 -908 2283 -904
rect 2256 -924 2260 -908
rect 2112 -945 2138 -941
rect 2147 -945 2151 -924
rect 2241 -945 2245 -934
rect 2147 -949 2245 -945
rect 523 -965 527 -949
rect 508 -1002 512 -975
rect -209 -1006 512 -1002
rect 1252 -1021 1256 -949
rect 1299 -994 1303 -949
rect 1402 -965 1406 -949
rect 1387 -994 1391 -975
rect 1299 -998 1391 -994
rect -209 -1025 1256 -1021
rect 2013 -1038 2017 -949
rect 2067 -994 2071 -949
rect 2170 -965 2174 -949
rect 2155 -994 2159 -975
rect 2067 -998 2159 -994
rect -209 -1042 2017 -1038
rect 127 -1096 327 -1092
rect 62 -1112 139 -1108
rect -183 -1144 17 -1140
rect -248 -1160 -171 -1156
rect -248 -1227 -244 -1160
rect -175 -1183 -171 -1160
rect -152 -1162 -148 -1144
rect -119 -1162 -115 -1144
rect -175 -1187 -151 -1183
rect -142 -1187 -138 -1166
rect -142 -1191 -74 -1187
rect -225 -1195 -188 -1191
rect -225 -1210 -221 -1195
rect -192 -1210 -188 -1195
rect -119 -1207 -115 -1191
rect -243 -1232 -224 -1228
rect -248 -1401 -244 -1232
rect -215 -1235 -211 -1214
rect -134 -1235 -130 -1217
rect -215 -1239 -130 -1235
rect -192 -1255 -188 -1239
rect -207 -1292 -203 -1265
rect -223 -1296 -203 -1292
rect -162 -1292 -158 -1239
rect -144 -1253 -96 -1249
rect -78 -1251 -74 -1191
rect -51 -1230 -47 -1144
rect -18 -1230 -14 -1144
rect -137 -1271 -133 -1253
rect -104 -1271 -100 -1253
rect -78 -1255 -50 -1251
rect -41 -1257 -37 -1234
rect -41 -1261 2 -1257
rect -18 -1275 -14 -1261
rect -162 -1296 -136 -1292
rect -127 -1296 -123 -1275
rect -33 -1296 -29 -1285
rect -207 -1345 -203 -1296
rect -127 -1300 -29 -1296
rect -104 -1316 -100 -1300
rect -119 -1345 -115 -1326
rect -207 -1351 -115 -1345
rect 13 -1358 17 -1144
rect 62 -1183 66 -1112
rect 135 -1135 139 -1112
rect 158 -1114 162 -1096
rect 191 -1114 195 -1096
rect 135 -1139 159 -1135
rect 168 -1139 172 -1118
rect 168 -1143 236 -1139
rect 85 -1147 122 -1143
rect 85 -1162 89 -1147
rect 118 -1162 122 -1147
rect 191 -1159 195 -1143
rect 37 -1187 86 -1183
rect 95 -1187 99 -1166
rect 176 -1187 180 -1169
rect 62 -1350 66 -1187
rect 95 -1191 180 -1187
rect 118 -1207 122 -1191
rect 103 -1244 107 -1217
rect 87 -1248 107 -1244
rect 148 -1244 152 -1191
rect 166 -1205 214 -1201
rect 232 -1203 236 -1143
rect 259 -1182 263 -1096
rect 292 -1182 296 -1096
rect 323 -1143 327 -1096
rect 870 -1099 1070 -1095
rect 1629 -1099 1829 -1095
rect 2365 -1099 2565 -1095
rect 805 -1115 882 -1111
rect 323 -1147 555 -1143
rect 560 -1147 760 -1143
rect 173 -1223 177 -1205
rect 206 -1223 210 -1205
rect 232 -1207 260 -1203
rect 269 -1207 273 -1186
rect 269 -1211 312 -1207
rect 292 -1227 296 -1211
rect 148 -1248 174 -1244
rect 183 -1248 187 -1227
rect 277 -1248 281 -1237
rect 103 -1297 107 -1248
rect 183 -1252 281 -1248
rect 206 -1268 210 -1252
rect 191 -1297 195 -1278
rect 103 -1301 195 -1297
rect 323 -1307 327 -1147
rect 495 -1163 572 -1159
rect 495 -1234 499 -1163
rect 568 -1186 572 -1163
rect 591 -1165 595 -1147
rect 624 -1165 628 -1147
rect 568 -1190 592 -1186
rect 601 -1190 605 -1169
rect 601 -1194 669 -1190
rect 518 -1198 555 -1194
rect 518 -1213 522 -1198
rect 551 -1213 555 -1198
rect 624 -1210 628 -1194
rect 452 -1238 519 -1234
rect 528 -1238 532 -1217
rect 609 -1238 613 -1220
rect 145 -1311 376 -1307
rect 145 -1329 149 -1311
rect 178 -1329 182 -1311
rect 211 -1329 215 -1311
rect 304 -1329 308 -1311
rect 372 -1329 376 -1311
rect 62 -1354 146 -1350
rect 155 -1354 159 -1333
rect 221 -1351 225 -1333
rect 155 -1358 212 -1354
rect 221 -1355 305 -1351
rect -166 -1362 17 -1358
rect -166 -1380 -162 -1362
rect -133 -1380 -129 -1362
rect -100 -1380 -96 -1362
rect 128 -1366 167 -1362
rect 178 -1374 182 -1358
rect 221 -1374 225 -1355
rect 301 -1363 326 -1359
rect 339 -1367 343 -1333
rect 382 -1354 386 -1333
rect 452 -1354 456 -1238
rect 382 -1358 456 -1354
rect 314 -1371 373 -1367
rect 314 -1377 318 -1371
rect 382 -1377 386 -1358
rect -248 -1405 -165 -1401
rect -156 -1405 -152 -1384
rect -156 -1409 -99 -1405
rect -182 -1417 -144 -1413
rect -133 -1425 -129 -1409
rect -90 -1410 -86 -1384
rect 145 -1393 149 -1378
rect 211 -1393 215 -1378
rect 304 -1393 308 -1381
rect 337 -1393 341 -1381
rect 372 -1393 376 -1381
rect 138 -1397 376 -1393
rect -90 -1414 237 -1410
rect -90 -1425 -86 -1414
rect -166 -1441 -162 -1429
rect -100 -1441 -96 -1429
rect -166 -1445 -96 -1441
rect 372 -1444 376 -1397
rect 495 -1404 499 -1238
rect 528 -1242 613 -1238
rect 551 -1258 555 -1242
rect 536 -1295 540 -1268
rect 520 -1299 540 -1295
rect 581 -1295 585 -1242
rect 599 -1256 647 -1252
rect 665 -1254 669 -1194
rect 692 -1233 696 -1147
rect 725 -1233 729 -1147
rect 606 -1274 610 -1256
rect 639 -1274 643 -1256
rect 665 -1258 693 -1254
rect 702 -1260 706 -1237
rect 702 -1264 745 -1260
rect 725 -1278 729 -1264
rect 581 -1299 607 -1295
rect 616 -1299 620 -1278
rect 710 -1299 714 -1288
rect 536 -1348 540 -1299
rect 616 -1303 714 -1299
rect 639 -1319 643 -1303
rect 624 -1348 628 -1329
rect 536 -1352 628 -1348
rect 756 -1361 760 -1147
rect 805 -1186 809 -1115
rect 878 -1138 882 -1115
rect 901 -1117 905 -1099
rect 934 -1117 938 -1099
rect 878 -1142 902 -1138
rect 911 -1142 915 -1121
rect 911 -1146 979 -1142
rect 828 -1150 865 -1146
rect 828 -1165 832 -1150
rect 861 -1165 865 -1150
rect 934 -1162 938 -1146
rect 780 -1190 829 -1186
rect 838 -1190 842 -1169
rect 919 -1190 923 -1172
rect 805 -1353 809 -1190
rect 838 -1194 923 -1190
rect 861 -1210 865 -1194
rect 846 -1247 850 -1220
rect 830 -1251 850 -1247
rect 891 -1247 895 -1194
rect 909 -1208 957 -1204
rect 975 -1206 979 -1146
rect 1002 -1185 1006 -1099
rect 1035 -1185 1039 -1099
rect 1066 -1143 1070 -1099
rect 1564 -1115 1641 -1111
rect 1066 -1147 1314 -1143
rect 1319 -1147 1519 -1143
rect 916 -1226 920 -1208
rect 949 -1226 953 -1208
rect 975 -1210 1003 -1206
rect 1012 -1210 1016 -1189
rect 1012 -1214 1055 -1210
rect 1035 -1230 1039 -1214
rect 891 -1251 917 -1247
rect 926 -1251 930 -1230
rect 1020 -1251 1024 -1240
rect 846 -1300 850 -1251
rect 926 -1255 1024 -1251
rect 949 -1271 953 -1255
rect 934 -1300 938 -1281
rect 846 -1304 938 -1300
rect 1066 -1310 1070 -1147
rect 1254 -1163 1331 -1159
rect 1254 -1234 1258 -1163
rect 1327 -1186 1331 -1163
rect 1350 -1165 1354 -1147
rect 1383 -1165 1387 -1147
rect 1327 -1190 1351 -1186
rect 1360 -1190 1364 -1169
rect 1360 -1194 1428 -1190
rect 1277 -1198 1314 -1194
rect 1277 -1213 1281 -1198
rect 1310 -1213 1314 -1198
rect 1383 -1210 1387 -1194
rect 1205 -1238 1278 -1234
rect 1287 -1238 1291 -1217
rect 1368 -1238 1372 -1220
rect 888 -1314 1119 -1310
rect 888 -1332 892 -1314
rect 921 -1332 925 -1314
rect 954 -1332 958 -1314
rect 1047 -1332 1051 -1314
rect 1115 -1332 1119 -1314
rect 805 -1357 889 -1353
rect 898 -1357 902 -1336
rect 964 -1354 968 -1336
rect 898 -1361 955 -1357
rect 964 -1358 1048 -1354
rect 577 -1365 760 -1361
rect 577 -1383 581 -1365
rect 610 -1383 614 -1365
rect 643 -1383 647 -1365
rect 871 -1369 910 -1365
rect 921 -1377 925 -1361
rect 964 -1377 968 -1358
rect 1044 -1366 1069 -1362
rect 1082 -1370 1086 -1336
rect 1125 -1357 1129 -1336
rect 1205 -1357 1209 -1238
rect 1125 -1361 1209 -1357
rect 1057 -1374 1116 -1370
rect 1057 -1380 1061 -1374
rect 1125 -1380 1129 -1361
rect 495 -1408 578 -1404
rect 587 -1408 591 -1387
rect 587 -1412 644 -1408
rect 561 -1420 599 -1416
rect 610 -1428 614 -1412
rect 653 -1413 657 -1387
rect 888 -1396 892 -1381
rect 954 -1396 958 -1381
rect 1047 -1396 1051 -1384
rect 1080 -1396 1084 -1384
rect 1115 -1396 1119 -1384
rect 881 -1400 1119 -1396
rect 653 -1417 980 -1413
rect 653 -1428 657 -1417
rect 577 -1444 581 -1432
rect 643 -1444 647 -1432
rect 1115 -1443 1119 -1400
rect 1254 -1404 1258 -1238
rect 1287 -1242 1372 -1238
rect 1310 -1258 1314 -1242
rect 1295 -1295 1299 -1268
rect 1279 -1299 1299 -1295
rect 1340 -1295 1344 -1242
rect 1358 -1256 1406 -1252
rect 1424 -1254 1428 -1194
rect 1451 -1233 1455 -1147
rect 1484 -1233 1488 -1147
rect 1365 -1274 1369 -1256
rect 1398 -1274 1402 -1256
rect 1424 -1258 1452 -1254
rect 1461 -1260 1465 -1237
rect 1461 -1264 1504 -1260
rect 1484 -1278 1488 -1264
rect 1340 -1299 1366 -1295
rect 1375 -1299 1379 -1278
rect 1469 -1299 1473 -1288
rect 1295 -1348 1299 -1299
rect 1375 -1303 1473 -1299
rect 1398 -1319 1402 -1303
rect 1383 -1348 1387 -1329
rect 1295 -1352 1387 -1348
rect 1299 -1354 1387 -1352
rect 1515 -1361 1519 -1147
rect 1564 -1186 1568 -1115
rect 1637 -1138 1641 -1115
rect 1660 -1117 1664 -1099
rect 1693 -1117 1697 -1099
rect 1637 -1142 1661 -1138
rect 1670 -1142 1674 -1121
rect 1670 -1146 1738 -1142
rect 1587 -1150 1624 -1146
rect 1587 -1165 1591 -1150
rect 1620 -1165 1624 -1150
rect 1693 -1162 1697 -1146
rect 1564 -1190 1588 -1186
rect 1597 -1190 1601 -1169
rect 1678 -1190 1682 -1172
rect 1564 -1353 1568 -1190
rect 1597 -1194 1682 -1190
rect 1620 -1210 1624 -1194
rect 1605 -1247 1609 -1220
rect 1589 -1251 1609 -1247
rect 1650 -1247 1654 -1194
rect 1668 -1208 1716 -1204
rect 1734 -1206 1738 -1146
rect 1761 -1185 1765 -1099
rect 1794 -1185 1798 -1099
rect 1825 -1143 1829 -1099
rect 2300 -1115 2377 -1111
rect 1825 -1147 2050 -1143
rect 2055 -1147 2255 -1143
rect 1675 -1226 1679 -1208
rect 1708 -1226 1712 -1208
rect 1734 -1210 1762 -1206
rect 1771 -1210 1775 -1189
rect 1771 -1214 1814 -1210
rect 1794 -1230 1798 -1214
rect 1650 -1251 1676 -1247
rect 1685 -1251 1689 -1230
rect 1779 -1251 1783 -1240
rect 1605 -1300 1609 -1251
rect 1685 -1255 1783 -1251
rect 1708 -1271 1712 -1255
rect 1825 -1277 1829 -1147
rect 1990 -1163 2067 -1159
rect 1990 -1234 1994 -1163
rect 2063 -1186 2067 -1163
rect 2086 -1165 2090 -1147
rect 2119 -1165 2123 -1147
rect 2063 -1190 2087 -1186
rect 2096 -1190 2100 -1169
rect 2096 -1194 2164 -1190
rect 2013 -1198 2050 -1194
rect 2013 -1213 2017 -1198
rect 2046 -1213 2050 -1198
rect 2119 -1210 2123 -1194
rect 1799 -1281 1829 -1277
rect 1935 -1238 2014 -1234
rect 2023 -1238 2027 -1217
rect 2104 -1238 2108 -1220
rect 1693 -1300 1697 -1281
rect 1605 -1304 1697 -1300
rect 1799 -1310 1803 -1281
rect 1647 -1314 1878 -1310
rect 1647 -1332 1651 -1314
rect 1680 -1332 1684 -1314
rect 1713 -1332 1717 -1314
rect 1806 -1332 1810 -1314
rect 1874 -1332 1878 -1314
rect 1564 -1357 1648 -1353
rect 1657 -1357 1661 -1336
rect 1723 -1354 1727 -1336
rect 1657 -1361 1714 -1357
rect 1723 -1358 1807 -1354
rect 1336 -1365 1519 -1361
rect 1336 -1383 1340 -1365
rect 1369 -1383 1373 -1365
rect 1402 -1383 1406 -1365
rect 1630 -1369 1669 -1365
rect 1680 -1377 1684 -1361
rect 1723 -1377 1727 -1358
rect 1803 -1366 1828 -1362
rect 1841 -1370 1845 -1336
rect 1884 -1357 1888 -1336
rect 1935 -1357 1939 -1238
rect 1884 -1361 1939 -1357
rect 1816 -1374 1875 -1370
rect 1816 -1380 1820 -1374
rect 1884 -1380 1888 -1361
rect 1254 -1408 1337 -1404
rect 1346 -1408 1350 -1387
rect 1346 -1412 1403 -1408
rect 1320 -1420 1358 -1416
rect 1369 -1428 1373 -1412
rect 1412 -1413 1416 -1387
rect 1647 -1396 1651 -1381
rect 1713 -1396 1717 -1381
rect 1806 -1396 1810 -1384
rect 1839 -1396 1843 -1384
rect 1874 -1396 1878 -1384
rect 1640 -1400 1878 -1396
rect 1412 -1417 1739 -1413
rect 1412 -1428 1416 -1417
rect 1336 -1443 1340 -1432
rect 1402 -1442 1406 -1432
rect 372 -1448 647 -1444
rect 1115 -1447 1401 -1443
rect 1874 -1443 1878 -1400
rect 1990 -1404 1994 -1238
rect 2023 -1242 2108 -1238
rect 2046 -1258 2050 -1242
rect 2031 -1295 2035 -1268
rect 2015 -1299 2035 -1295
rect 2076 -1295 2080 -1242
rect 2094 -1256 2142 -1252
rect 2160 -1254 2164 -1194
rect 2187 -1233 2191 -1147
rect 2220 -1233 2224 -1147
rect 2101 -1274 2105 -1256
rect 2134 -1274 2138 -1256
rect 2160 -1258 2188 -1254
rect 2197 -1260 2201 -1237
rect 2197 -1264 2240 -1260
rect 2220 -1278 2224 -1264
rect 2076 -1299 2102 -1295
rect 2111 -1299 2115 -1278
rect 2205 -1299 2209 -1288
rect 2031 -1348 2035 -1299
rect 2111 -1303 2209 -1299
rect 2134 -1319 2138 -1303
rect 2119 -1348 2123 -1329
rect 2031 -1352 2123 -1348
rect 2035 -1354 2123 -1352
rect 2251 -1361 2255 -1147
rect 2300 -1186 2304 -1115
rect 2373 -1138 2377 -1115
rect 2396 -1117 2400 -1099
rect 2429 -1117 2433 -1099
rect 2373 -1142 2397 -1138
rect 2406 -1142 2410 -1121
rect 2406 -1146 2474 -1142
rect 2323 -1150 2360 -1146
rect 2323 -1165 2327 -1150
rect 2356 -1165 2360 -1150
rect 2429 -1162 2433 -1146
rect 2300 -1190 2324 -1186
rect 2333 -1190 2337 -1169
rect 2414 -1190 2418 -1172
rect 2300 -1353 2304 -1190
rect 2333 -1194 2418 -1190
rect 2356 -1210 2360 -1194
rect 2341 -1247 2345 -1220
rect 2325 -1251 2345 -1247
rect 2386 -1247 2390 -1194
rect 2404 -1208 2452 -1204
rect 2470 -1206 2474 -1146
rect 2497 -1185 2501 -1099
rect 2530 -1185 2534 -1099
rect 2411 -1226 2415 -1208
rect 2444 -1226 2448 -1208
rect 2470 -1210 2498 -1206
rect 2507 -1210 2511 -1189
rect 2507 -1214 2550 -1210
rect 2530 -1230 2534 -1214
rect 2386 -1251 2412 -1247
rect 2421 -1251 2425 -1230
rect 2515 -1251 2519 -1240
rect 2341 -1300 2345 -1251
rect 2421 -1255 2519 -1251
rect 2444 -1271 2448 -1255
rect 2561 -1277 2565 -1099
rect 2535 -1281 2565 -1277
rect 2429 -1300 2433 -1281
rect 2341 -1304 2433 -1300
rect 2535 -1310 2539 -1281
rect 2383 -1314 2614 -1310
rect 2383 -1332 2387 -1314
rect 2416 -1332 2420 -1314
rect 2449 -1332 2453 -1314
rect 2542 -1332 2546 -1314
rect 2610 -1332 2614 -1314
rect 2300 -1357 2384 -1353
rect 2393 -1357 2397 -1336
rect 2459 -1354 2463 -1336
rect 2393 -1361 2450 -1357
rect 2459 -1358 2543 -1354
rect 2072 -1365 2255 -1361
rect 2072 -1383 2076 -1365
rect 2105 -1383 2109 -1365
rect 2138 -1383 2142 -1365
rect 2366 -1369 2405 -1365
rect 2416 -1377 2420 -1361
rect 2459 -1377 2463 -1358
rect 2539 -1366 2564 -1362
rect 2577 -1370 2581 -1336
rect 2620 -1357 2624 -1336
rect 2620 -1361 2632 -1357
rect 2552 -1374 2611 -1370
rect 2552 -1380 2556 -1374
rect 2620 -1380 2624 -1361
rect 1990 -1408 2073 -1404
rect 2082 -1408 2086 -1387
rect 2082 -1412 2139 -1408
rect 2056 -1420 2094 -1416
rect 2105 -1428 2109 -1412
rect 2148 -1413 2152 -1387
rect 2383 -1396 2387 -1381
rect 2449 -1396 2453 -1381
rect 2542 -1396 2546 -1384
rect 2575 -1396 2579 -1384
rect 2610 -1396 2614 -1384
rect 2376 -1400 2614 -1396
rect 2148 -1417 2475 -1413
rect 2148 -1428 2152 -1417
rect 2072 -1443 2076 -1432
rect 2138 -1441 2142 -1432
rect 1874 -1446 2137 -1443
rect -245 -1463 467 -1459
rect 1241 -1476 1245 -1472
rect -245 -1480 1245 -1476
rect 1965 -1488 1969 -1483
rect -245 -1492 1969 -1488
rect -504 -1589 -388 -1585
rect -504 -1600 -500 -1589
rect -580 -1614 -576 -1604
rect -514 -1614 -510 -1604
rect -580 -1618 -510 -1614
rect -450 -1642 -250 -1638
rect -234 -1642 1180 -1638
rect -608 -1708 -604 -1644
rect -588 -1657 -60 -1653
rect -579 -1675 -575 -1657
rect -546 -1675 -542 -1657
rect -513 -1675 -509 -1657
rect -461 -1667 -218 -1663
rect -202 -1667 787 -1663
rect -588 -1700 -578 -1696
rect -569 -1700 -565 -1679
rect -569 -1704 -512 -1700
rect -608 -1712 -557 -1708
rect -608 -1800 -604 -1712
rect -546 -1720 -542 -1704
rect -503 -1705 -499 -1679
rect -472 -1692 -186 -1688
rect -170 -1692 415 -1688
rect -503 -1709 -151 -1705
rect -135 -1709 -125 -1705
rect -503 -1720 -499 -1709
rect -579 -1734 -575 -1724
rect -513 -1734 -509 -1724
rect -579 -1738 -509 -1734
rect -588 -1748 -512 -1744
rect -582 -1767 -578 -1748
rect -549 -1767 -545 -1748
rect -516 -1767 -512 -1748
rect -588 -1792 -581 -1788
rect -572 -1792 -568 -1771
rect -572 -1796 -515 -1792
rect -608 -1804 -560 -1800
rect -608 -1892 -604 -1804
rect -549 -1812 -545 -1796
rect -506 -1797 -502 -1771
rect -506 -1801 -473 -1797
rect -129 -1800 -125 -1709
rect -17 -1713 152 -1709
rect -78 -1729 -5 -1725
rect -78 -1800 -74 -1729
rect -9 -1752 -5 -1729
rect 14 -1731 18 -1713
rect 47 -1731 51 -1713
rect -9 -1756 15 -1752
rect 24 -1756 28 -1735
rect 24 -1760 92 -1756
rect -59 -1764 -22 -1760
rect -59 -1779 -55 -1764
rect -26 -1779 -22 -1764
rect 47 -1776 51 -1760
rect -506 -1812 -502 -1801
rect -129 -1804 -58 -1800
rect -49 -1804 -45 -1783
rect 32 -1804 36 -1786
rect -49 -1808 36 -1804
rect -582 -1826 -578 -1816
rect -516 -1826 -512 -1816
rect -26 -1824 -22 -1808
rect -582 -1830 -512 -1826
rect -588 -1840 -512 -1836
rect -582 -1859 -578 -1840
rect -549 -1859 -545 -1840
rect -516 -1859 -512 -1840
rect -477 -1846 -101 -1842
rect -588 -1884 -581 -1880
rect -572 -1884 -568 -1863
rect -572 -1888 -515 -1884
rect -608 -1896 -560 -1892
rect -608 -1984 -604 -1896
rect -549 -1904 -545 -1888
rect -506 -1889 -502 -1863
rect -506 -1893 -462 -1889
rect -506 -1904 -502 -1893
rect -41 -1896 -37 -1834
rect 4 -1861 8 -1808
rect 29 -1822 70 -1818
rect 88 -1820 92 -1760
rect 115 -1799 119 -1713
rect 148 -1781 152 -1713
rect 407 -1725 415 -1692
rect 472 -1713 641 -1709
rect 407 -1729 484 -1725
rect 148 -1785 245 -1781
rect 148 -1799 152 -1785
rect 241 -1803 245 -1785
rect 407 -1800 415 -1729
rect 480 -1752 484 -1729
rect 503 -1731 507 -1713
rect 536 -1731 540 -1713
rect 480 -1756 504 -1752
rect 513 -1756 517 -1735
rect 513 -1760 581 -1756
rect 430 -1764 467 -1760
rect 430 -1779 434 -1764
rect 463 -1779 467 -1764
rect 536 -1776 540 -1760
rect 29 -1840 33 -1822
rect 62 -1840 66 -1822
rect 88 -1824 116 -1820
rect 125 -1824 129 -1803
rect 125 -1828 242 -1824
rect 251 -1828 255 -1807
rect 407 -1808 431 -1800
rect 440 -1804 444 -1783
rect 521 -1804 525 -1786
rect 440 -1808 525 -1804
rect 463 -1824 467 -1808
rect 148 -1844 152 -1828
rect 251 -1832 287 -1828
rect 251 -1842 255 -1832
rect 4 -1865 30 -1861
rect 39 -1865 43 -1844
rect 133 -1865 137 -1854
rect 39 -1869 137 -1865
rect 62 -1885 66 -1869
rect 241 -1879 245 -1846
rect 448 -1861 452 -1834
rect 128 -1883 245 -1879
rect 407 -1869 452 -1861
rect 493 -1861 497 -1808
rect 511 -1822 559 -1818
rect 577 -1820 581 -1760
rect 604 -1799 608 -1713
rect 637 -1781 641 -1713
rect 637 -1785 681 -1781
rect 637 -1799 641 -1785
rect 677 -1803 681 -1785
rect 779 -1800 787 -1667
rect 856 -1713 1059 -1709
rect 795 -1729 868 -1725
rect 795 -1800 799 -1729
rect 864 -1752 868 -1729
rect 887 -1731 891 -1713
rect 920 -1731 924 -1713
rect 864 -1756 888 -1752
rect 897 -1756 901 -1735
rect 897 -1760 965 -1756
rect 814 -1764 851 -1760
rect 814 -1779 818 -1764
rect 847 -1779 851 -1764
rect 920 -1776 924 -1760
rect 518 -1840 522 -1822
rect 551 -1840 555 -1822
rect 577 -1824 605 -1820
rect 614 -1824 618 -1803
rect 614 -1828 678 -1824
rect 687 -1828 691 -1807
rect 779 -1808 815 -1800
rect 824 -1804 828 -1783
rect 905 -1804 909 -1786
rect 824 -1808 909 -1804
rect 847 -1824 851 -1808
rect 637 -1844 641 -1828
rect 687 -1832 703 -1828
rect 687 -1842 691 -1832
rect 493 -1865 519 -1861
rect 528 -1865 532 -1844
rect 622 -1865 626 -1854
rect 528 -1869 626 -1865
rect -388 -1904 -119 -1896
rect -103 -1904 -37 -1896
rect -582 -1918 -578 -1908
rect -516 -1918 -512 -1908
rect -582 -1922 -512 -1918
rect -588 -1932 -512 -1928
rect -582 -1951 -578 -1932
rect -549 -1951 -545 -1932
rect -516 -1951 -512 -1932
rect -588 -1976 -581 -1972
rect -572 -1976 -568 -1955
rect -572 -1980 -515 -1976
rect -608 -1988 -560 -1984
rect -608 -2075 -604 -1988
rect -549 -1996 -545 -1980
rect -506 -1981 -502 -1955
rect -506 -1985 -494 -1981
rect -506 -1996 -502 -1985
rect -498 -1991 -494 -1985
rect -456 -1991 -451 -1990
rect -498 -1995 -451 -1991
rect -582 -2010 -578 -2000
rect -516 -2010 -512 -2000
rect -582 -2014 -512 -2010
rect -586 -2024 -507 -2020
rect -577 -2042 -573 -2024
rect -544 -2042 -540 -2024
rect -511 -2042 -507 -2024
rect -586 -2067 -576 -2063
rect -567 -2067 -563 -2046
rect -567 -2071 -510 -2067
rect -608 -2079 -555 -2075
rect -608 -2167 -604 -2079
rect -544 -2087 -540 -2071
rect -501 -2072 -497 -2046
rect -388 -2072 -384 -1904
rect -41 -1914 -37 -1904
rect 47 -1914 51 -1895
rect -41 -1918 51 -1914
rect 98 -1913 102 -1890
rect 407 -1924 415 -1869
rect 448 -1914 452 -1869
rect 551 -1885 555 -1869
rect 677 -1879 681 -1846
rect 832 -1861 836 -1834
rect 617 -1883 681 -1879
rect 812 -1869 836 -1861
rect 877 -1861 881 -1808
rect 895 -1822 943 -1818
rect 961 -1820 965 -1760
rect 1022 -1799 1026 -1713
rect 1055 -1781 1059 -1713
rect 1055 -1785 1099 -1781
rect 1055 -1799 1059 -1785
rect 1095 -1803 1099 -1785
rect 902 -1840 906 -1822
rect 935 -1840 939 -1822
rect 961 -1824 1023 -1820
rect 1032 -1824 1036 -1803
rect 1032 -1828 1096 -1824
rect 1105 -1828 1109 -1807
rect 1176 -1824 1180 -1642
rect 1271 -1737 1440 -1733
rect 1210 -1753 1283 -1749
rect 1210 -1824 1214 -1753
rect 1279 -1776 1283 -1753
rect 1302 -1755 1306 -1737
rect 1335 -1755 1339 -1737
rect 1279 -1780 1303 -1776
rect 1312 -1780 1316 -1759
rect 1312 -1784 1380 -1780
rect 1229 -1788 1266 -1784
rect 1229 -1803 1233 -1788
rect 1262 -1803 1266 -1788
rect 1335 -1800 1339 -1784
rect 1055 -1844 1059 -1828
rect 1105 -1832 1153 -1828
rect 1176 -1828 1230 -1824
rect 1239 -1828 1243 -1807
rect 1320 -1828 1324 -1810
rect 1239 -1832 1324 -1828
rect 1105 -1842 1109 -1832
rect 877 -1865 903 -1861
rect 912 -1865 916 -1844
rect 1040 -1865 1044 -1854
rect 912 -1869 1044 -1865
rect 536 -1914 540 -1895
rect 448 -1918 540 -1914
rect -501 -2076 -384 -2072
rect -340 -1932 209 -1924
rect 225 -1932 415 -1924
rect -501 -2087 -497 -2076
rect -577 -2101 -573 -2091
rect -511 -2101 -507 -2091
rect -577 -2105 -507 -2101
rect -586 -2115 -510 -2111
rect -580 -2134 -576 -2115
rect -547 -2134 -543 -2115
rect -514 -2134 -510 -2115
rect -586 -2159 -579 -2155
rect -570 -2159 -566 -2138
rect -570 -2163 -513 -2159
rect -608 -2171 -558 -2167
rect -608 -2259 -604 -2171
rect -547 -2179 -543 -2163
rect -504 -2164 -500 -2138
rect -340 -2164 -336 -1932
rect 812 -1952 820 -1869
rect 832 -1914 836 -1869
rect 935 -1885 939 -1869
rect 1095 -1879 1099 -1846
rect 1262 -1848 1266 -1832
rect 1035 -1883 1099 -1879
rect 1247 -1885 1251 -1858
rect 1168 -1889 1251 -1885
rect 1292 -1885 1296 -1832
rect 1317 -1846 1358 -1842
rect 1376 -1844 1380 -1784
rect 1403 -1823 1407 -1737
rect 1436 -1801 1440 -1737
rect 1436 -1805 1475 -1801
rect 1436 -1823 1440 -1805
rect 1471 -1823 1475 -1805
rect 1317 -1864 1321 -1846
rect 1350 -1864 1354 -1846
rect 1376 -1848 1404 -1844
rect 1413 -1848 1417 -1827
rect 1481 -1848 1485 -1827
rect 1413 -1852 1472 -1848
rect 1481 -1852 1493 -1848
rect 1436 -1868 1440 -1852
rect 1481 -1862 1485 -1852
rect 1292 -1889 1318 -1885
rect 1327 -1889 1331 -1868
rect 1471 -1876 1475 -1866
rect 1421 -1889 1425 -1878
rect 1464 -1880 1475 -1876
rect 920 -1914 924 -1895
rect 832 -1918 924 -1914
rect -504 -2168 -336 -2164
rect -316 -1960 624 -1952
rect 640 -1960 820 -1952
rect -504 -2179 -500 -2168
rect -580 -2193 -576 -2183
rect -514 -2193 -510 -2183
rect -580 -2197 -510 -2193
rect -586 -2207 -510 -2203
rect -580 -2226 -576 -2207
rect -547 -2226 -543 -2207
rect -514 -2226 -510 -2207
rect -586 -2251 -579 -2247
rect -570 -2251 -566 -2230
rect -570 -2255 -513 -2251
rect -608 -2263 -558 -2259
rect -608 -2351 -604 -2263
rect -547 -2271 -543 -2255
rect -504 -2259 -500 -2230
rect -316 -2259 -312 -1960
rect 1168 -1980 1176 -1889
rect 1247 -1938 1251 -1889
rect 1327 -1893 1425 -1889
rect 1350 -1909 1354 -1893
rect 1335 -1938 1339 -1919
rect 1247 -1942 1339 -1938
rect -504 -2263 -312 -2259
rect -268 -1983 1176 -1980
rect -268 -1988 1068 -1983
rect 1073 -1988 1176 -1983
rect -504 -2271 -500 -2263
rect -580 -2285 -576 -2275
rect -514 -2285 -510 -2275
rect -580 -2289 -510 -2285
rect -586 -2299 -510 -2295
rect -580 -2318 -576 -2299
rect -547 -2318 -543 -2299
rect -514 -2318 -510 -2299
rect -586 -2343 -579 -2339
rect -570 -2343 -566 -2322
rect -570 -2347 -513 -2343
rect -608 -2355 -558 -2351
rect -547 -2363 -543 -2347
rect -504 -2348 -500 -2322
rect -268 -2348 -264 -1988
rect -165 -2004 199 -1996
rect -197 -2021 618 -2013
rect 612 -2024 618 -2021
rect -208 -2046 1062 -2038
rect 1056 -2049 1062 -2046
rect 120 -2071 842 -2067
rect 847 -2071 1435 -2067
rect -67 -2138 31 -2130
rect -67 -2158 -59 -2138
rect -135 -2166 -59 -2158
rect -67 -2187 -59 -2166
rect -33 -2148 3 -2144
rect -33 -2166 -29 -2148
rect -1 -2151 3 -2148
rect -67 -2191 -32 -2187
rect -23 -2191 -19 -2170
rect -5 -2173 -1 -2152
rect -5 -2177 23 -2173
rect -23 -2195 11 -2191
rect -23 -2205 -19 -2195
rect -33 -2219 -29 -2209
rect -48 -2223 -29 -2219
rect -52 -2312 -48 -2223
rect -35 -2234 -12 -2230
rect -35 -2259 -31 -2234
rect -25 -2284 -21 -2263
rect -38 -2288 -34 -2284
rect -25 -2288 -13 -2284
rect -25 -2298 -21 -2288
rect -35 -2312 -31 -2302
rect 7 -2311 11 -2195
rect 19 -2256 23 -2177
rect 27 -2208 31 -2138
rect 120 -2152 124 -2071
rect 47 -2156 124 -2152
rect 54 -2174 58 -2156
rect 87 -2174 91 -2156
rect 120 -2174 124 -2156
rect 199 -2107 205 -2084
rect 334 -2089 338 -2071
rect 389 -2089 393 -2071
rect 442 -2089 446 -2071
rect 477 -2084 481 -2071
rect 199 -2111 335 -2107
rect 199 -2167 205 -2111
rect 247 -2128 260 -2124
rect 256 -2142 260 -2128
rect 199 -2171 257 -2167
rect 266 -2172 270 -2146
rect 348 -2143 352 -2093
rect 407 -2143 411 -2093
rect 452 -2131 456 -2093
rect 452 -2135 512 -2131
rect 348 -2147 443 -2143
rect 407 -2163 411 -2147
rect 452 -2163 456 -2135
rect 51 -2199 55 -2195
rect 64 -2199 68 -2178
rect 64 -2203 121 -2199
rect 27 -2212 44 -2208
rect 40 -2241 44 -2212
rect 87 -2219 91 -2203
rect 130 -2204 134 -2178
rect 266 -2176 321 -2172
rect 266 -2187 270 -2176
rect 130 -2208 167 -2204
rect 256 -2204 260 -2191
rect 317 -2193 321 -2176
rect 334 -2177 338 -2167
rect 442 -2177 446 -2167
rect 334 -2181 450 -2177
rect 334 -2204 338 -2181
rect 477 -2204 481 -2167
rect 200 -2208 338 -2204
rect 352 -2208 481 -2204
rect 130 -2219 134 -2208
rect 72 -2241 76 -2229
rect 40 -2245 76 -2241
rect 19 -2260 125 -2256
rect 55 -2290 59 -2260
rect 88 -2290 92 -2260
rect 121 -2290 125 -2260
rect -52 -2316 -6 -2312
rect 7 -2315 56 -2311
rect 65 -2315 69 -2294
rect -504 -2352 -264 -2348
rect -504 -2363 -500 -2352
rect -12 -2356 -6 -2316
rect 65 -2319 122 -2315
rect 41 -2357 45 -2324
rect 88 -2335 92 -2319
rect 131 -2320 135 -2294
rect 131 -2324 150 -2320
rect 131 -2335 135 -2324
rect 73 -2357 77 -2345
rect 41 -2361 77 -2357
rect -580 -2377 -576 -2367
rect -514 -2377 -510 -2367
rect -580 -2381 -510 -2377
rect 159 -2380 167 -2208
rect 238 -2220 260 -2216
rect 234 -2326 238 -2220
rect 256 -2234 260 -2220
rect 253 -2266 257 -2262
rect 266 -2279 270 -2238
rect 256 -2293 260 -2283
rect 281 -2293 285 -2208
rect 317 -2244 321 -2217
rect 352 -2226 356 -2208
rect 407 -2226 411 -2208
rect 460 -2226 464 -2208
rect 317 -2248 353 -2244
rect 366 -2280 370 -2230
rect 425 -2280 429 -2230
rect 470 -2268 474 -2230
rect 470 -2272 498 -2268
rect 366 -2284 461 -2280
rect 256 -2298 285 -2293
rect 425 -2300 429 -2284
rect 470 -2300 474 -2272
rect 352 -2314 356 -2304
rect 460 -2314 464 -2304
rect 352 -2318 464 -2314
rect -42 -2388 167 -2380
rect 204 -2330 238 -2326
rect 204 -2384 215 -2330
rect -42 -2510 -34 -2388
rect 508 -2396 512 -2135
rect 541 -2289 545 -2071
rect 612 -2107 618 -2084
rect 750 -2089 754 -2071
rect 805 -2089 809 -2071
rect 858 -2089 862 -2071
rect 612 -2111 751 -2107
rect 612 -2167 618 -2111
rect 663 -2128 676 -2124
rect 672 -2142 676 -2128
rect 612 -2171 673 -2167
rect 682 -2172 686 -2146
rect 764 -2143 768 -2093
rect 823 -2143 827 -2093
rect 868 -2131 872 -2093
rect 868 -2135 916 -2131
rect 764 -2147 859 -2143
rect 823 -2163 827 -2147
rect 868 -2163 872 -2135
rect 682 -2176 737 -2172
rect 682 -2187 686 -2176
rect 672 -2232 676 -2191
rect 733 -2193 737 -2176
rect 750 -2177 754 -2167
rect 858 -2177 862 -2167
rect 750 -2181 862 -2177
rect 750 -2232 754 -2181
rect 858 -2208 862 -2181
rect 613 -2236 754 -2232
rect 768 -2224 843 -2220
rect 654 -2248 669 -2244
rect 665 -2262 669 -2248
rect 541 -2293 618 -2289
rect 548 -2311 552 -2293
rect 581 -2311 585 -2293
rect 614 -2311 618 -2293
rect 662 -2294 666 -2290
rect 675 -2307 679 -2266
rect 524 -2336 549 -2332
rect 558 -2336 562 -2315
rect 538 -2369 542 -2336
rect 558 -2340 615 -2336
rect 550 -2348 570 -2344
rect 581 -2356 585 -2340
rect 624 -2341 628 -2315
rect 665 -2322 669 -2311
rect 697 -2322 701 -2236
rect 733 -2272 737 -2245
rect 768 -2254 772 -2224
rect 823 -2254 827 -2224
rect 848 -2224 880 -2220
rect 876 -2254 880 -2224
rect 733 -2276 769 -2272
rect 782 -2308 786 -2258
rect 841 -2308 845 -2258
rect 886 -2296 890 -2258
rect 886 -2300 898 -2296
rect 782 -2312 877 -2308
rect 665 -2326 756 -2322
rect 624 -2345 663 -2341
rect 624 -2356 628 -2345
rect 548 -2368 552 -2360
rect 614 -2368 618 -2360
rect 681 -2368 685 -2326
rect 752 -2342 756 -2326
rect 841 -2328 845 -2312
rect 886 -2328 890 -2300
rect 768 -2342 772 -2332
rect 876 -2342 880 -2332
rect 752 -2346 880 -2342
rect 548 -2372 685 -2368
rect -26 -2404 512 -2396
rect -26 -2502 -18 -2404
rect 908 -2412 916 -2135
rect 950 -2250 954 -2071
rect 1056 -2107 1062 -2084
rect 1200 -2089 1204 -2071
rect 1255 -2089 1259 -2071
rect 1308 -2072 1435 -2071
rect 1308 -2089 1312 -2072
rect 1056 -2111 1201 -2107
rect 1056 -2167 1062 -2111
rect 1107 -2128 1120 -2124
rect 1116 -2142 1120 -2128
rect 1056 -2171 1117 -2167
rect 1126 -2172 1130 -2146
rect 1214 -2143 1218 -2093
rect 1273 -2143 1277 -2093
rect 1318 -2131 1322 -2093
rect 1318 -2135 1366 -2131
rect 1214 -2147 1309 -2143
rect 1273 -2163 1277 -2147
rect 1318 -2163 1322 -2135
rect 1126 -2176 1187 -2172
rect 1126 -2187 1130 -2176
rect 1116 -2204 1120 -2191
rect 1183 -2193 1187 -2176
rect 1200 -2177 1204 -2167
rect 1308 -2177 1312 -2167
rect 1200 -2181 1312 -2177
rect 1200 -2204 1204 -2181
rect 1057 -2208 1204 -2204
rect 1218 -2208 1330 -2204
rect 950 -2254 1027 -2250
rect 957 -2272 961 -2254
rect 990 -2272 994 -2254
rect 1023 -2272 1027 -2254
rect 942 -2297 958 -2293
rect 967 -2297 971 -2276
rect 943 -2323 947 -2297
rect 967 -2301 1024 -2297
rect 959 -2309 979 -2305
rect 990 -2317 994 -2301
rect 1033 -2302 1037 -2276
rect 1033 -2306 1052 -2302
rect 1033 -2317 1037 -2306
rect 957 -2331 961 -2321
rect 1023 -2331 1027 -2321
rect 957 -2335 1027 -2331
rect 1048 -2340 1052 -2306
rect 1058 -2314 1062 -2208
rect 1098 -2220 1119 -2216
rect 1115 -2234 1119 -2220
rect 1112 -2263 1116 -2259
rect 1125 -2279 1129 -2238
rect 1115 -2295 1119 -2283
rect 1141 -2295 1145 -2208
rect 1183 -2244 1187 -2217
rect 1218 -2226 1222 -2208
rect 1273 -2226 1277 -2208
rect 1326 -2226 1330 -2208
rect 1183 -2248 1219 -2244
rect 1232 -2280 1236 -2230
rect 1291 -2280 1295 -2230
rect 1336 -2268 1340 -2230
rect 1336 -2272 1348 -2268
rect 1232 -2284 1327 -2280
rect 1115 -2299 1145 -2295
rect 1291 -2300 1295 -2284
rect 1336 -2300 1340 -2272
rect 1218 -2314 1222 -2304
rect 1326 -2314 1330 -2304
rect 1058 -2318 1330 -2314
rect 1058 -2330 1062 -2318
rect -10 -2420 916 -2412
rect -10 -2494 -2 -2420
rect 1358 -2428 1366 -2135
rect 1431 -2245 1435 -2072
rect 1431 -2249 1566 -2245
rect 1438 -2267 1442 -2249
rect 1489 -2267 1493 -2249
rect 1530 -2267 1534 -2249
rect 1562 -2267 1566 -2249
rect 1435 -2289 1439 -2285
rect 1448 -2293 1452 -2271
rect 1509 -2285 1513 -2271
rect 1509 -2289 1534 -2285
rect 1530 -2293 1534 -2289
rect 1448 -2297 1563 -2293
rect 1435 -2305 1468 -2301
rect 1435 -2314 1492 -2310
rect 1435 -2323 1516 -2319
rect 1530 -2329 1534 -2297
rect 1572 -2310 1576 -2271
rect 1572 -2314 1584 -2310
rect 1572 -2329 1576 -2314
rect 1438 -2341 1442 -2333
rect 1562 -2341 1566 -2333
rect 1389 -2345 1566 -2341
rect 6 -2436 1366 -2428
rect 6 -2486 14 -2436
rect 36 -2450 441 -2446
rect 36 -2468 40 -2450
rect 167 -2468 171 -2450
rect 306 -2468 310 -2450
rect 437 -2468 441 -2450
rect 6 -2490 37 -2486
rect -10 -2498 58 -2494
rect -26 -2506 79 -2502
rect -42 -2514 100 -2510
rect 120 -2518 124 -2472
rect 177 -2489 181 -2472
rect 177 -2493 189 -2489
rect 297 -2490 307 -2486
rect 46 -2522 168 -2518
rect 46 -2536 50 -2522
rect 120 -2526 124 -2522
rect 93 -2530 124 -2526
rect 93 -2536 97 -2530
rect 177 -2536 181 -2493
rect 297 -2499 328 -2495
rect 297 -2508 349 -2504
rect 297 -2517 370 -2513
rect 390 -2521 394 -2472
rect 447 -2503 451 -2472
rect 447 -2508 458 -2503
rect 316 -2525 438 -2521
rect 316 -2539 320 -2525
rect 390 -2529 394 -2525
rect 363 -2533 394 -2529
rect 363 -2539 367 -2533
rect 447 -2539 451 -2508
rect 36 -2553 40 -2540
rect 69 -2553 73 -2540
rect 167 -2553 171 -2540
rect 306 -2553 310 -2543
rect 339 -2553 343 -2543
rect 437 -2553 441 -2543
rect 9 -2556 441 -2553
rect -608 -2635 -604 -2571
rect -588 -2584 -77 -2580
rect -579 -2602 -575 -2584
rect -546 -2602 -542 -2584
rect -513 -2602 -509 -2584
rect -588 -2627 -578 -2623
rect -569 -2627 -565 -2606
rect -569 -2631 -512 -2627
rect -608 -2639 -557 -2635
rect -608 -2727 -604 -2639
rect -546 -2647 -542 -2631
rect -503 -2632 -499 -2606
rect -503 -2636 -94 -2632
rect -503 -2647 -499 -2636
rect -579 -2661 -575 -2651
rect -513 -2661 -509 -2651
rect -579 -2665 -509 -2661
rect -588 -2675 -512 -2671
rect -582 -2694 -578 -2675
rect -549 -2694 -545 -2675
rect -516 -2694 -512 -2675
rect -588 -2719 -581 -2715
rect -572 -2719 -568 -2698
rect -572 -2723 -515 -2719
rect -608 -2731 -560 -2727
rect -608 -2819 -604 -2731
rect -549 -2739 -545 -2723
rect -506 -2724 -502 -2698
rect -506 -2728 -107 -2724
rect -506 -2739 -502 -2728
rect -582 -2753 -578 -2743
rect -516 -2753 -512 -2743
rect -582 -2757 -512 -2753
rect -588 -2767 -512 -2763
rect -582 -2786 -578 -2767
rect -549 -2786 -545 -2767
rect -516 -2786 -512 -2767
rect -588 -2811 -581 -2807
rect -572 -2811 -568 -2790
rect -572 -2815 -515 -2811
rect -608 -2823 -560 -2819
rect -608 -2911 -604 -2823
rect -549 -2831 -545 -2815
rect -506 -2816 -502 -2790
rect -506 -2820 -133 -2816
rect -506 -2831 -502 -2820
rect -582 -2845 -578 -2835
rect -516 -2845 -512 -2835
rect -582 -2849 -512 -2845
rect -588 -2859 -512 -2855
rect -582 -2878 -578 -2859
rect -549 -2878 -545 -2859
rect -516 -2878 -512 -2859
rect -588 -2903 -581 -2899
rect -572 -2903 -568 -2882
rect -572 -2907 -515 -2903
rect -608 -2915 -560 -2911
rect -608 -3002 -604 -2915
rect -549 -2923 -545 -2907
rect -506 -2908 -502 -2882
rect -506 -2912 -161 -2908
rect -506 -2923 -502 -2912
rect -582 -2937 -578 -2927
rect -516 -2937 -512 -2927
rect -582 -2941 -512 -2937
rect -586 -2951 -507 -2947
rect -577 -2969 -573 -2951
rect -544 -2969 -540 -2951
rect -511 -2969 -507 -2951
rect -586 -2994 -576 -2990
rect -567 -2994 -563 -2973
rect -567 -2998 -510 -2994
rect -608 -3006 -555 -3002
rect -608 -3094 -604 -3006
rect -544 -3014 -540 -2998
rect -501 -2999 -497 -2973
rect -501 -3003 -477 -2999
rect -501 -3014 -497 -3003
rect -577 -3028 -573 -3018
rect -511 -3028 -507 -3018
rect -577 -3032 -507 -3028
rect -586 -3042 -510 -3038
rect -580 -3061 -576 -3042
rect -547 -3061 -543 -3042
rect -514 -3061 -510 -3042
rect -165 -3060 -161 -2912
rect -137 -2967 -133 -2820
rect -111 -2875 -107 -2728
rect -98 -2782 -94 -2636
rect -81 -2739 -77 -2584
rect -81 -2743 26 -2739
rect -81 -2761 -77 -2743
rect -48 -2761 -44 -2743
rect -15 -2761 -11 -2743
rect -98 -2786 -80 -2782
rect -71 -2786 -67 -2765
rect -71 -2790 -14 -2786
rect -86 -2798 -59 -2794
rect -48 -2806 -44 -2790
rect -5 -2791 -1 -2765
rect -5 -2795 6 -2791
rect -5 -2806 -1 -2795
rect -81 -2820 -77 -2810
rect -15 -2820 -11 -2810
rect -81 -2824 -11 -2820
rect 22 -2832 26 -2743
rect -81 -2836 26 -2832
rect -81 -2854 -77 -2836
rect -48 -2854 -44 -2836
rect -15 -2854 -11 -2836
rect -111 -2879 -80 -2875
rect -71 -2879 -67 -2858
rect -71 -2883 -14 -2879
rect -86 -2891 -59 -2887
rect -48 -2899 -44 -2883
rect -5 -2884 -1 -2858
rect -5 -2888 6 -2884
rect -5 -2899 -1 -2888
rect -81 -2913 -77 -2903
rect -15 -2913 -11 -2903
rect -81 -2917 -11 -2913
rect 22 -2924 26 -2836
rect -81 -2928 26 -2924
rect -81 -2946 -77 -2928
rect -48 -2946 -44 -2928
rect -15 -2946 -11 -2928
rect -137 -2971 -80 -2967
rect -71 -2971 -67 -2950
rect -71 -2975 -14 -2971
rect -86 -2983 -59 -2979
rect -48 -2991 -44 -2975
rect -5 -2976 -1 -2950
rect -5 -2980 6 -2976
rect -5 -2991 -1 -2980
rect -81 -3005 -77 -2995
rect -15 -3005 -11 -2995
rect -81 -3009 -11 -3005
rect 22 -3017 26 -2928
rect -81 -3021 26 -3017
rect -81 -3039 -77 -3021
rect -48 -3039 -44 -3021
rect -15 -3039 -11 -3021
rect -165 -3064 -80 -3060
rect -71 -3064 -67 -3043
rect -586 -3086 -579 -3082
rect -570 -3086 -566 -3065
rect -570 -3090 -513 -3086
rect -608 -3098 -558 -3094
rect -608 -3186 -604 -3098
rect -547 -3106 -543 -3090
rect -504 -3091 -500 -3065
rect -71 -3068 -14 -3064
rect -86 -3076 -59 -3072
rect -48 -3084 -44 -3068
rect -5 -3069 -1 -3043
rect -5 -3073 6 -3069
rect -5 -3084 -1 -3073
rect -504 -3095 -477 -3091
rect -504 -3106 -500 -3095
rect -81 -3098 -77 -3088
rect -15 -3098 -11 -3088
rect -81 -3102 -11 -3098
rect -580 -3120 -576 -3110
rect -514 -3120 -510 -3110
rect -580 -3124 -510 -3120
rect -586 -3134 -510 -3130
rect -580 -3153 -576 -3134
rect -547 -3153 -543 -3134
rect -514 -3153 -510 -3134
rect -586 -3178 -579 -3174
rect -570 -3178 -566 -3157
rect -570 -3182 -513 -3178
rect -608 -3190 -558 -3186
rect -608 -3278 -604 -3190
rect -547 -3198 -543 -3182
rect -504 -3186 -500 -3157
rect -504 -3190 -477 -3186
rect -504 -3198 -500 -3190
rect -580 -3212 -576 -3202
rect -514 -3212 -510 -3202
rect -580 -3216 -510 -3212
rect -586 -3226 -510 -3222
rect -580 -3245 -576 -3226
rect -547 -3245 -543 -3226
rect -514 -3245 -510 -3226
rect -586 -3270 -579 -3266
rect -570 -3270 -566 -3249
rect -570 -3274 -513 -3270
rect -608 -3282 -558 -3278
rect -547 -3290 -543 -3274
rect -504 -3275 -500 -3249
rect -504 -3279 -477 -3275
rect -504 -3290 -500 -3279
rect -580 -3304 -576 -3294
rect -514 -3304 -510 -3294
rect -580 -3308 -510 -3304
<< m2contact >>
rect -809 120 -804 125
rect -821 62 -816 67
rect -893 11 -888 16
rect -829 11 -824 16
rect -846 6 -841 11
rect -820 -1 -815 4
rect -942 -89 -937 -84
rect -639 120 -634 125
rect -643 11 -638 16
rect -449 11 -444 16
rect -423 11 -418 16
rect -548 2 -543 7
rect -691 -61 -686 -56
rect -915 -1643 -910 -1638
rect -937 -2570 -932 -2565
rect -884 -787 -879 -782
rect -884 -1580 -879 -1575
rect -884 -2343 -879 -2338
rect -864 -695 -859 -690
rect -864 -1488 -859 -1483
rect -864 -2251 -859 -2246
rect -844 -603 -839 -598
rect -844 -1396 -839 -1391
rect -844 -2159 -839 -2154
rect -824 -511 -819 -506
rect -824 -1304 -819 -1299
rect -824 -2067 -819 -2062
rect -804 -420 -799 -415
rect -804 -1213 -799 -1208
rect -804 -1976 -799 -1971
rect -784 -328 -779 -323
rect -784 -1121 -779 -1116
rect -784 -1884 -779 -1879
rect -764 -236 -759 -231
rect -764 -1029 -759 -1024
rect -764 -1792 -759 -1787
rect -744 -144 -739 -139
rect -487 -90 -482 -85
rect -593 -144 -588 -139
rect -330 -129 -325 -124
rect -188 0 -183 5
rect 410 0 415 5
rect 1289 0 1294 5
rect 2057 0 2062 5
rect -257 -91 -248 -86
rect -193 -47 -188 -42
rect -153 -72 -148 -67
rect -226 -120 -221 -115
rect -307 -148 -302 -142
rect -478 -153 -473 -148
rect -96 -109 -91 -104
rect -56 -66 -51 -61
rect 341 -91 350 -86
rect 405 -47 410 -42
rect 445 -72 450 -67
rect 372 -120 377 -115
rect -52 -140 -47 -135
rect 502 -109 507 -104
rect 542 -66 547 -61
rect 1220 -91 1229 -86
rect 1284 -47 1289 -42
rect 1324 -72 1329 -67
rect 1251 -120 1256 -115
rect 546 -140 551 -135
rect -509 -182 -504 -177
rect -138 -181 -133 -176
rect -593 -236 -588 -231
rect -469 -245 -464 -240
rect -512 -274 -507 -269
rect -593 -328 -588 -323
rect -461 -337 -456 -332
rect -512 -366 -507 -361
rect -593 -420 -588 -415
rect -512 -458 -507 -453
rect -591 -511 -586 -506
rect -507 -549 -502 -544
rect -591 -603 -586 -598
rect -510 -641 -505 -636
rect -591 -695 -586 -690
rect -510 -733 -505 -728
rect -591 -787 -586 -782
rect 1381 -109 1386 -104
rect 1421 -66 1426 -61
rect 1988 -91 1997 -86
rect 2052 -47 2057 -42
rect 2092 -72 2097 -67
rect 2019 -120 2024 -115
rect 1425 -140 1430 -135
rect 2149 -109 2154 -104
rect 2189 -66 2194 -61
rect 2193 -140 2198 -135
rect 460 -181 465 -176
rect 1339 -181 1344 -176
rect 2107 -181 2112 -176
rect 93 -303 98 -298
rect -217 -351 -212 -346
rect -222 -398 -217 -393
rect -182 -423 -177 -418
rect -255 -471 -250 -466
rect -125 -460 -120 -455
rect -85 -417 -80 -412
rect -27 -468 -22 -463
rect -81 -491 -76 -486
rect -252 -508 -247 -503
rect -167 -532 -162 -527
rect 88 -350 93 -345
rect 128 -375 133 -370
rect 55 -423 60 -418
rect 185 -412 190 -407
rect 225 -369 230 -364
rect 836 -306 841 -301
rect 1595 -306 1600 -301
rect 2331 -306 2336 -301
rect 526 -354 531 -349
rect 283 -418 288 -413
rect 229 -443 234 -438
rect 58 -460 63 -455
rect 143 -484 148 -479
rect 521 -401 526 -396
rect 561 -426 566 -421
rect 94 -574 99 -569
rect -216 -625 -211 -620
rect 110 -610 115 -604
rect 208 -621 213 -616
rect -125 -652 -120 -647
rect 488 -474 493 -469
rect 618 -463 623 -458
rect 658 -420 663 -415
rect 716 -471 721 -466
rect 662 -494 667 -489
rect 491 -511 496 -506
rect 576 -535 581 -530
rect 831 -353 836 -348
rect 871 -378 876 -373
rect 798 -426 803 -421
rect 928 -415 933 -410
rect 968 -372 973 -367
rect 1285 -354 1290 -349
rect 1026 -421 1031 -416
rect 972 -446 977 -441
rect 801 -463 806 -458
rect 886 -487 891 -482
rect 1280 -401 1285 -396
rect 1320 -426 1325 -421
rect 837 -577 842 -572
rect 527 -628 532 -623
rect 853 -613 858 -607
rect 951 -624 956 -619
rect 1247 -474 1252 -469
rect 1377 -463 1382 -458
rect 1417 -420 1422 -415
rect 1475 -471 1480 -466
rect 1421 -494 1426 -489
rect 1250 -511 1255 -506
rect 1335 -535 1340 -530
rect 1590 -353 1595 -348
rect 1630 -378 1635 -373
rect 1557 -426 1562 -421
rect 1687 -415 1692 -410
rect 1727 -372 1732 -367
rect 2021 -354 2026 -349
rect 1785 -421 1790 -416
rect 1731 -446 1736 -441
rect 1560 -463 1565 -458
rect 1645 -487 1650 -482
rect 2016 -401 2021 -396
rect 2056 -426 2061 -421
rect 1596 -577 1601 -572
rect 1286 -628 1291 -623
rect 1612 -613 1617 -607
rect 1710 -624 1715 -619
rect 618 -655 623 -650
rect 1372 -654 1377 -649
rect 1983 -474 1988 -469
rect 2113 -463 2118 -458
rect 2153 -420 2158 -415
rect 2211 -471 2216 -466
rect 2157 -494 2162 -489
rect 1986 -511 1991 -506
rect 2071 -535 2076 -530
rect 2326 -353 2331 -348
rect 2366 -378 2371 -373
rect 2293 -426 2298 -421
rect 2423 -415 2428 -410
rect 2463 -372 2468 -367
rect 2521 -421 2526 -416
rect 2467 -446 2472 -441
rect 2296 -463 2301 -458
rect 2381 -487 2386 -482
rect 2332 -577 2337 -572
rect 2022 -628 2027 -623
rect 2348 -613 2353 -607
rect 2446 -624 2451 -619
rect 2108 -653 2113 -648
rect -279 -670 -274 -665
rect 438 -670 443 -665
rect 1211 -679 1216 -674
rect -279 -687 -274 -682
rect 1936 -690 1941 -685
rect -279 -699 -274 -694
rect -337 -808 -332 -803
rect -510 -825 -505 -820
rect -744 -937 -739 -932
rect -159 -793 -154 -788
rect 439 -793 444 -788
rect 1318 -793 1323 -788
rect 2086 -793 2091 -788
rect -228 -884 -219 -879
rect -164 -840 -159 -835
rect -124 -865 -119 -860
rect -593 -937 -588 -932
rect -404 -922 -399 -917
rect -321 -922 -316 -917
rect -197 -913 -192 -908
rect -278 -941 -273 -935
rect -478 -946 -473 -941
rect -67 -902 -62 -897
rect -27 -859 -22 -854
rect 370 -884 379 -879
rect 434 -840 439 -835
rect 474 -865 479 -860
rect 401 -913 406 -908
rect -23 -933 -18 -928
rect 531 -902 536 -897
rect 571 -859 576 -854
rect 1249 -884 1258 -879
rect 1313 -840 1318 -835
rect 1353 -865 1358 -860
rect 1280 -913 1285 -908
rect 575 -933 580 -928
rect -509 -975 -504 -970
rect -109 -974 -104 -969
rect -593 -1029 -588 -1024
rect -469 -1038 -464 -1033
rect -512 -1067 -507 -1062
rect -593 -1121 -588 -1116
rect -461 -1130 -456 -1125
rect -512 -1159 -507 -1154
rect -593 -1213 -588 -1208
rect -512 -1251 -507 -1246
rect -591 -1304 -586 -1299
rect -507 -1342 -502 -1337
rect -591 -1396 -586 -1391
rect -510 -1434 -505 -1429
rect -591 -1488 -586 -1483
rect -510 -1526 -505 -1521
rect -591 -1580 -586 -1575
rect 1410 -902 1415 -897
rect 1450 -859 1455 -854
rect 2017 -884 2026 -879
rect 2081 -840 2086 -835
rect 2121 -865 2126 -860
rect 2048 -913 2053 -908
rect 1454 -933 1459 -928
rect 2178 -902 2183 -897
rect 2218 -859 2223 -854
rect 2222 -933 2227 -928
rect 489 -974 494 -969
rect 1368 -974 1373 -969
rect 2136 -974 2141 -969
rect 122 -1096 127 -1091
rect -188 -1144 -183 -1139
rect -193 -1191 -188 -1186
rect -153 -1216 -148 -1211
rect -226 -1264 -221 -1259
rect -96 -1253 -91 -1248
rect -56 -1210 -51 -1205
rect 2 -1261 7 -1256
rect -52 -1284 -47 -1279
rect -223 -1301 -218 -1296
rect -138 -1325 -133 -1320
rect 117 -1143 122 -1138
rect 157 -1168 162 -1163
rect 84 -1216 89 -1211
rect 214 -1205 219 -1200
rect 254 -1162 259 -1157
rect 865 -1099 870 -1094
rect 1624 -1099 1629 -1094
rect 2360 -1099 2365 -1094
rect 555 -1147 560 -1142
rect 312 -1211 317 -1206
rect 258 -1236 263 -1231
rect 87 -1253 92 -1248
rect 172 -1277 177 -1272
rect 550 -1194 555 -1189
rect 590 -1219 595 -1214
rect 123 -1367 128 -1362
rect -187 -1418 -182 -1413
rect 139 -1403 144 -1397
rect 237 -1414 242 -1409
rect -96 -1445 -91 -1440
rect 517 -1267 522 -1262
rect 647 -1256 652 -1251
rect 687 -1213 692 -1208
rect 745 -1264 750 -1259
rect 691 -1287 696 -1282
rect 520 -1304 525 -1299
rect 605 -1328 610 -1323
rect 860 -1146 865 -1141
rect 900 -1171 905 -1166
rect 827 -1219 832 -1214
rect 957 -1208 962 -1203
rect 997 -1165 1002 -1160
rect 1314 -1147 1319 -1142
rect 1055 -1214 1060 -1209
rect 1001 -1239 1006 -1234
rect 830 -1256 835 -1251
rect 915 -1280 920 -1275
rect 1309 -1194 1314 -1189
rect 1349 -1219 1354 -1214
rect 866 -1370 871 -1365
rect 556 -1421 561 -1416
rect 882 -1406 887 -1400
rect 980 -1417 985 -1412
rect 1276 -1267 1281 -1262
rect 1406 -1256 1411 -1251
rect 1446 -1213 1451 -1208
rect 1504 -1264 1509 -1259
rect 1450 -1287 1455 -1282
rect 1279 -1304 1284 -1299
rect 1364 -1328 1369 -1323
rect 1619 -1146 1624 -1141
rect 1659 -1171 1664 -1166
rect 1586 -1219 1591 -1214
rect 1716 -1208 1721 -1203
rect 1756 -1165 1761 -1160
rect 2050 -1147 2055 -1142
rect 1814 -1214 1819 -1209
rect 1760 -1239 1765 -1234
rect 1589 -1256 1594 -1251
rect 1674 -1280 1679 -1275
rect 2045 -1194 2050 -1189
rect 2085 -1219 2090 -1214
rect 1625 -1370 1630 -1365
rect 1315 -1421 1320 -1416
rect 1641 -1406 1646 -1400
rect 1739 -1417 1744 -1412
rect 647 -1448 652 -1443
rect 1401 -1447 1406 -1442
rect 2012 -1267 2017 -1262
rect 2142 -1256 2147 -1251
rect 2182 -1213 2187 -1208
rect 2240 -1264 2245 -1259
rect 2186 -1287 2191 -1282
rect 2015 -1304 2020 -1299
rect 2100 -1328 2105 -1323
rect 2355 -1146 2360 -1141
rect 2395 -1171 2400 -1166
rect 2322 -1219 2327 -1214
rect 2452 -1208 2457 -1203
rect 2492 -1165 2497 -1160
rect 2550 -1214 2555 -1209
rect 2496 -1239 2501 -1234
rect 2325 -1256 2330 -1251
rect 2410 -1280 2415 -1275
rect 2361 -1370 2366 -1365
rect 2051 -1421 2056 -1416
rect 2377 -1406 2382 -1400
rect 2475 -1417 2480 -1412
rect 2137 -1446 2142 -1441
rect -250 -1463 -245 -1458
rect 467 -1463 472 -1458
rect 1240 -1472 1245 -1467
rect -250 -1480 -245 -1475
rect 1965 -1483 1970 -1478
rect -250 -1492 -245 -1487
rect -510 -1618 -505 -1613
rect -455 -1642 -450 -1637
rect -250 -1642 -234 -1637
rect -744 -1700 -739 -1695
rect -604 -1648 -599 -1643
rect -60 -1657 -55 -1652
rect -466 -1667 -461 -1662
rect -218 -1667 -202 -1662
rect -593 -1700 -588 -1695
rect -477 -1692 -472 -1687
rect -186 -1692 -170 -1687
rect -151 -1709 -135 -1704
rect -509 -1738 -504 -1733
rect -593 -1792 -588 -1787
rect -478 -1797 -473 -1792
rect -22 -1713 -17 -1708
rect -27 -1760 -22 -1755
rect 13 -1785 18 -1780
rect -512 -1830 -507 -1825
rect -60 -1833 -55 -1828
rect -482 -1846 -477 -1841
rect -101 -1846 -96 -1841
rect -593 -1884 -588 -1879
rect -467 -1889 -462 -1884
rect 70 -1822 75 -1817
rect 110 -1779 115 -1774
rect 467 -1713 472 -1708
rect 462 -1760 467 -1755
rect 502 -1785 507 -1780
rect 429 -1833 434 -1828
rect 114 -1853 119 -1848
rect 123 -1883 128 -1878
rect 559 -1822 564 -1817
rect 599 -1779 604 -1774
rect 851 -1713 856 -1708
rect 846 -1760 851 -1755
rect 886 -1785 891 -1780
rect 813 -1833 818 -1828
rect 603 -1853 608 -1848
rect 28 -1894 33 -1889
rect 98 -1890 103 -1885
rect -119 -1904 -103 -1896
rect -512 -1922 -507 -1917
rect -593 -1976 -588 -1971
rect -456 -1990 -451 -1985
rect -512 -2014 -507 -2009
rect -591 -2067 -586 -2062
rect 98 -1918 106 -1913
rect 612 -1883 617 -1878
rect 943 -1822 948 -1817
rect 1017 -1779 1022 -1774
rect 1266 -1737 1271 -1732
rect 1261 -1784 1266 -1779
rect 1301 -1809 1306 -1804
rect 1021 -1853 1026 -1848
rect 517 -1894 522 -1889
rect 209 -1932 225 -1924
rect -507 -2105 -502 -2100
rect -591 -2159 -586 -2154
rect 1030 -1883 1035 -1878
rect 1228 -1857 1233 -1852
rect 1358 -1846 1363 -1841
rect 1398 -1803 1403 -1798
rect 1402 -1877 1407 -1872
rect 1464 -1885 1469 -1880
rect 901 -1894 906 -1889
rect 624 -1960 640 -1952
rect -510 -2197 -505 -2192
rect -591 -2251 -586 -2246
rect 1316 -1918 1321 -1913
rect 1068 -1988 1073 -1983
rect -510 -2289 -505 -2284
rect -591 -2343 -586 -2338
rect -170 -2004 -165 -1996
rect 199 -2005 205 -1996
rect -202 -2021 -197 -2013
rect 612 -2033 618 -2024
rect -213 -2046 -208 -2038
rect 1056 -2058 1062 -2049
rect 842 -2071 847 -2066
rect -151 -2166 -135 -2158
rect -1 -2156 4 -2151
rect -53 -2223 -48 -2218
rect -12 -2234 -7 -2229
rect -43 -2288 -38 -2283
rect -13 -2288 -8 -2283
rect 42 -2156 47 -2151
rect 199 -2084 205 -2075
rect 242 -2076 247 -2071
rect 476 -2089 481 -2084
rect 242 -2128 247 -2123
rect 363 -2119 368 -2114
rect 476 -2167 481 -2162
rect 44 -2199 51 -2194
rect 195 -2208 200 -2203
rect 450 -2181 455 -2176
rect 317 -2198 322 -2193
rect 53 -2228 58 -2223
rect 119 -2228 124 -2223
rect 36 -2329 41 -2324
rect -6 -2356 -1 -2351
rect 150 -2324 155 -2319
rect 54 -2344 59 -2339
rect 120 -2344 125 -2339
rect -510 -2381 -505 -2376
rect 233 -2220 238 -2215
rect 248 -2266 253 -2261
rect 270 -2273 275 -2268
rect 317 -2217 322 -2212
rect 381 -2256 386 -2251
rect 498 -2272 503 -2267
rect 347 -2318 352 -2313
rect 204 -2389 215 -2384
rect 612 -2084 618 -2075
rect 658 -2076 663 -2071
rect 658 -2128 663 -2123
rect 779 -2119 784 -2114
rect 608 -2236 613 -2231
rect 733 -2198 738 -2193
rect 862 -2208 867 -2203
rect 649 -2248 654 -2243
rect 657 -2294 662 -2289
rect 679 -2288 684 -2283
rect 733 -2245 738 -2240
rect 843 -2225 848 -2220
rect 797 -2284 802 -2279
rect 898 -2300 903 -2295
rect 1056 -2084 1062 -2075
rect 1102 -2076 1107 -2071
rect 1291 -2076 1296 -2071
rect 1102 -2128 1107 -2123
rect 1229 -2119 1234 -2114
rect 1052 -2208 1057 -2203
rect 1183 -2198 1188 -2193
rect 1292 -2204 1297 -2199
rect 1027 -2335 1032 -2330
rect 1093 -2220 1098 -2215
rect 1107 -2263 1112 -2258
rect 1129 -2261 1134 -2256
rect 1183 -2217 1188 -2212
rect 1247 -2256 1252 -2251
rect 1348 -2272 1353 -2267
rect 1058 -2335 1063 -2330
rect 1388 -2341 1393 -2336
rect 204 -2446 215 -2441
rect 292 -2490 297 -2485
rect 292 -2499 297 -2494
rect 292 -2508 297 -2503
rect 292 -2517 297 -2512
rect 4 -2556 9 -2551
rect -744 -2627 -739 -2622
rect -604 -2575 -599 -2570
rect -593 -2627 -588 -2622
rect -764 -2719 -759 -2714
rect -509 -2665 -504 -2660
rect -593 -2719 -588 -2714
rect -784 -2811 -779 -2806
rect -512 -2757 -507 -2752
rect -593 -2811 -588 -2806
rect -804 -2903 -799 -2898
rect -512 -2849 -507 -2844
rect -593 -2903 -588 -2898
rect -824 -2994 -819 -2989
rect -512 -2941 -507 -2936
rect -591 -2994 -586 -2989
rect -844 -3086 -839 -3081
rect -477 -3003 -472 -2998
rect -507 -3032 -502 -3027
rect -91 -2798 -86 -2793
rect -11 -2824 -6 -2819
rect -91 -2891 -86 -2886
rect -11 -2917 -6 -2912
rect -91 -2983 -86 -2978
rect -11 -3009 -6 -3004
rect -591 -3086 -586 -3081
rect -864 -3178 -859 -3173
rect -91 -3076 -86 -3071
rect -477 -3095 -472 -3090
rect -11 -3102 -6 -3097
rect -510 -3124 -505 -3119
rect -591 -3178 -586 -3173
rect -884 -3270 -879 -3265
rect -477 -3190 -472 -3185
rect -510 -3216 -505 -3211
rect -591 -3270 -586 -3265
rect -477 -3279 -472 -3274
rect -510 -3308 -505 -3303
<< pdm12contact >>
rect 267 -570 272 -565
rect 1010 -573 1015 -568
rect 1769 -573 1774 -568
rect 2505 -573 2510 -568
rect 296 -1363 301 -1358
rect 1039 -1366 1044 -1361
rect 1798 -1366 1803 -1361
rect 2534 -1366 2539 -1361
<< metal2 >>
rect -837 175 -659 179
rect -837 124 -833 175
rect -837 120 -809 124
rect -663 124 -659 175
rect -663 120 -639 124
rect -897 -38 -893 15
rect -837 10 -833 120
rect -841 6 -833 10
rect -829 -38 -825 11
rect -820 4 -816 62
rect -666 11 -643 15
rect -485 11 -449 15
rect -361 15 1996 19
rect -418 11 -357 15
rect -666 -38 -662 11
rect -897 -42 -662 -38
rect -547 -47 -543 2
rect -941 -51 -543 -47
rect -941 -84 -937 -51
rect -485 -57 -481 11
rect -686 -61 -481 -57
rect -904 -73 -537 -69
rect -904 -884 -900 -73
rect -739 -144 -593 -140
rect -486 -178 -482 -90
rect -504 -182 -482 -178
rect -759 -236 -593 -232
rect -486 -270 -482 -182
rect -507 -274 -482 -270
rect -779 -328 -593 -324
rect -486 -362 -482 -274
rect -507 -366 -482 -362
rect -799 -420 -593 -416
rect -486 -454 -482 -366
rect -507 -458 -482 -454
rect -819 -511 -591 -507
rect -486 -545 -482 -458
rect -502 -549 -482 -545
rect -839 -603 -591 -599
rect -486 -637 -482 -549
rect -505 -641 -482 -637
rect -859 -695 -591 -691
rect -486 -729 -482 -641
rect -477 -695 -473 -153
rect -469 -683 -465 -245
rect -461 -666 -457 -337
rect -361 -512 -357 11
rect -257 -86 -253 15
rect -192 -42 -188 4
rect -91 -66 -56 -62
rect -225 -129 -221 -120
rect -152 -129 -148 -72
rect -91 -109 -87 -66
rect 341 -86 345 15
rect 406 -42 410 4
rect 507 -66 542 -62
rect 373 -129 377 -120
rect 446 -129 450 -72
rect 507 -109 511 -66
rect 1220 -86 1228 15
rect 1285 -42 1289 4
rect 1386 -66 1421 -62
rect 1252 -129 1256 -120
rect 1325 -129 1329 -72
rect 1386 -109 1390 -66
rect 1988 -86 1996 15
rect 2053 -42 2057 4
rect 2154 -66 2189 -62
rect 2020 -129 2024 -120
rect 2093 -129 2097 -72
rect 2154 -109 2158 -66
rect -350 -133 -148 -129
rect 366 -133 450 -129
rect 1245 -133 1329 -129
rect 2013 -133 2097 -129
rect -350 -480 -346 -133
rect -306 -299 -302 -148
rect -152 -190 -148 -133
rect -137 -190 -133 -181
rect -51 -190 -47 -140
rect 446 -190 450 -133
rect 461 -190 465 -181
rect 547 -190 551 -140
rect 1325 -190 1329 -133
rect 1340 -190 1344 -181
rect 1426 -190 1430 -140
rect 2093 -190 2097 -133
rect 2108 -190 2112 -181
rect 2194 -190 2198 -140
rect -152 -194 2198 -190
rect -306 -303 93 -299
rect -221 -393 -217 -303
rect 89 -345 93 -303
rect 522 -306 836 -302
rect 1281 -306 1595 -302
rect 2017 -306 2331 -302
rect 190 -369 225 -365
rect -120 -417 -85 -413
rect -254 -480 -250 -471
rect -181 -480 -177 -423
rect -120 -460 -116 -417
rect 56 -432 60 -423
rect 129 -432 133 -375
rect 190 -412 194 -369
rect 522 -396 526 -306
rect 832 -348 836 -306
rect 933 -372 968 -368
rect 288 -418 310 -414
rect 623 -420 658 -416
rect 56 -436 133 -432
rect 59 -464 63 -460
rect -22 -468 63 -464
rect -350 -484 -177 -480
rect -251 -512 -247 -508
rect -361 -516 -247 -512
rect -251 -620 -247 -516
rect -181 -541 -177 -484
rect -166 -541 -162 -532
rect -80 -541 -76 -491
rect -181 -545 -76 -541
rect -251 -624 -216 -620
rect -80 -648 -76 -545
rect 59 -569 63 -468
rect 129 -493 133 -436
rect 144 -493 148 -484
rect 230 -493 234 -443
rect 489 -483 493 -474
rect 562 -483 566 -426
rect 623 -463 627 -420
rect 799 -435 803 -426
rect 872 -435 876 -378
rect 933 -415 937 -372
rect 1281 -396 1285 -306
rect 1591 -348 1595 -306
rect 1692 -372 1727 -368
rect 1031 -421 1053 -417
rect 1382 -420 1417 -416
rect 799 -439 876 -435
rect 802 -467 806 -463
rect 721 -471 806 -467
rect 482 -487 566 -483
rect 129 -497 234 -493
rect 59 -573 94 -569
rect 230 -606 234 -497
rect 492 -515 496 -511
rect 443 -519 496 -515
rect 115 -610 234 -606
rect 242 -570 267 -566
rect 144 -648 148 -610
rect 242 -616 246 -570
rect 213 -620 246 -616
rect -120 -652 148 -648
rect -461 -670 -279 -666
rect 443 -670 447 -519
rect 492 -623 496 -519
rect 562 -544 566 -487
rect 577 -544 581 -535
rect 663 -544 667 -494
rect 562 -548 667 -544
rect 492 -627 527 -623
rect 663 -651 667 -548
rect 802 -572 806 -471
rect 872 -496 876 -439
rect 887 -496 891 -487
rect 973 -496 977 -446
rect 1248 -483 1252 -474
rect 1321 -483 1325 -426
rect 1382 -463 1386 -420
rect 1558 -435 1562 -426
rect 1631 -435 1635 -378
rect 1692 -415 1696 -372
rect 2017 -396 2021 -306
rect 2327 -348 2331 -306
rect 2428 -372 2463 -368
rect 1790 -421 1808 -417
rect 2118 -420 2153 -416
rect 1558 -439 1635 -435
rect 1561 -467 1565 -463
rect 1480 -471 1565 -467
rect 1248 -487 1325 -483
rect 872 -500 977 -496
rect 802 -576 837 -572
rect 973 -609 977 -500
rect 1251 -515 1255 -511
rect 1212 -519 1255 -515
rect 858 -613 977 -609
rect 985 -573 1010 -569
rect 887 -651 891 -613
rect 985 -619 989 -573
rect 956 -623 989 -619
rect 623 -655 891 -651
rect 1212 -674 1216 -519
rect 1251 -623 1255 -519
rect 1321 -544 1325 -487
rect 1336 -544 1340 -535
rect 1422 -544 1426 -494
rect 1321 -548 1426 -544
rect 1251 -627 1286 -623
rect 1422 -650 1426 -548
rect 1561 -572 1565 -471
rect 1631 -496 1635 -439
rect 1646 -496 1650 -487
rect 1732 -496 1736 -446
rect 1984 -483 1988 -474
rect 2057 -483 2061 -426
rect 2118 -463 2122 -420
rect 2294 -435 2298 -426
rect 2367 -435 2371 -378
rect 2428 -415 2432 -372
rect 2526 -421 2542 -417
rect 2294 -439 2371 -435
rect 2297 -467 2301 -463
rect 2216 -471 2301 -467
rect 1984 -487 2061 -483
rect 1631 -500 1736 -496
rect 1561 -576 1596 -572
rect 1732 -609 1736 -500
rect 1987 -515 1991 -511
rect 1936 -519 1991 -515
rect 1617 -613 1736 -609
rect 1744 -573 1769 -569
rect 1646 -650 1650 -613
rect 1744 -619 1748 -573
rect 1715 -623 1748 -619
rect 1377 -654 1650 -650
rect -469 -687 -279 -683
rect 1936 -685 1940 -519
rect 1987 -623 1991 -519
rect 2057 -544 2061 -487
rect 2072 -544 2076 -535
rect 2158 -544 2162 -494
rect 2057 -548 2162 -544
rect 1987 -627 2022 -623
rect 2158 -650 2162 -548
rect 2297 -572 2301 -471
rect 2367 -496 2371 -439
rect 2382 -496 2386 -487
rect 2468 -496 2472 -446
rect 2367 -500 2472 -496
rect 2297 -576 2332 -572
rect 2468 -609 2472 -500
rect 2353 -613 2472 -609
rect 2480 -573 2505 -569
rect 2382 -650 2386 -613
rect 2480 -619 2484 -573
rect 2451 -623 2484 -619
rect 2113 -653 2386 -650
rect -477 -699 -279 -695
rect -505 -733 -482 -729
rect -879 -787 -591 -783
rect -486 -821 -482 -733
rect -332 -778 2025 -774
rect -505 -825 -482 -821
rect -904 -888 -630 -884
rect -486 -918 -482 -825
rect -486 -922 -404 -918
rect -739 -937 -593 -933
rect -486 -971 -482 -922
rect -504 -975 -482 -971
rect -759 -1029 -593 -1025
rect -486 -1063 -482 -975
rect -507 -1067 -482 -1063
rect -779 -1121 -593 -1117
rect -486 -1155 -482 -1067
rect -507 -1159 -482 -1155
rect -799 -1213 -593 -1209
rect -486 -1247 -482 -1159
rect -507 -1251 -482 -1247
rect -819 -1304 -591 -1300
rect -486 -1338 -482 -1251
rect -502 -1342 -482 -1338
rect -839 -1396 -591 -1392
rect -486 -1430 -482 -1342
rect -505 -1434 -482 -1430
rect -859 -1488 -591 -1484
rect -486 -1522 -482 -1434
rect -477 -1488 -473 -946
rect -469 -1476 -465 -1038
rect -461 -1459 -457 -1130
rect -332 -1305 -328 -778
rect -228 -879 -224 -778
rect -163 -835 -159 -789
rect -62 -859 -27 -855
rect -196 -922 -192 -913
rect -123 -922 -119 -865
rect -62 -902 -58 -859
rect 370 -879 374 -778
rect 435 -835 439 -789
rect 536 -859 571 -855
rect 402 -922 406 -913
rect 475 -922 479 -865
rect 536 -902 540 -859
rect 1249 -879 1257 -778
rect 1314 -835 1318 -789
rect 1415 -859 1450 -855
rect 1281 -922 1285 -913
rect 1354 -922 1358 -865
rect 1415 -902 1419 -859
rect 2017 -879 2025 -778
rect 2082 -835 2086 -789
rect 2183 -859 2218 -855
rect 2049 -922 2053 -913
rect 2122 -922 2126 -865
rect 2183 -902 2187 -859
rect -321 -926 -119 -922
rect 395 -926 479 -922
rect 1274 -926 1358 -922
rect 2042 -926 2126 -922
rect -321 -1273 -317 -926
rect -277 -1092 -273 -941
rect -123 -983 -119 -926
rect -108 -983 -104 -974
rect -22 -983 -18 -933
rect 475 -983 479 -926
rect 490 -983 494 -974
rect 576 -983 580 -933
rect 1354 -983 1358 -926
rect 1369 -983 1373 -974
rect 1455 -983 1459 -933
rect 2122 -983 2126 -926
rect 2137 -983 2141 -974
rect 2223 -983 2227 -933
rect -123 -987 2227 -983
rect -277 -1096 122 -1092
rect -192 -1186 -188 -1096
rect 118 -1138 122 -1096
rect 551 -1099 865 -1095
rect 1310 -1099 1624 -1095
rect 2046 -1099 2360 -1095
rect 219 -1162 254 -1158
rect -91 -1210 -56 -1206
rect -225 -1273 -221 -1264
rect -152 -1273 -148 -1216
rect -91 -1253 -87 -1210
rect 85 -1225 89 -1216
rect 158 -1225 162 -1168
rect 219 -1205 223 -1162
rect 551 -1189 555 -1099
rect 861 -1141 865 -1099
rect 962 -1165 997 -1161
rect 317 -1211 339 -1207
rect 652 -1213 687 -1209
rect 85 -1229 162 -1225
rect 88 -1257 92 -1253
rect 7 -1261 92 -1257
rect -321 -1277 -148 -1273
rect -222 -1305 -218 -1301
rect -332 -1309 -218 -1305
rect -222 -1413 -218 -1309
rect -152 -1334 -148 -1277
rect -137 -1334 -133 -1325
rect -51 -1334 -47 -1284
rect -152 -1338 -47 -1334
rect -222 -1417 -187 -1413
rect -51 -1441 -47 -1338
rect 88 -1362 92 -1261
rect 158 -1286 162 -1229
rect 173 -1286 177 -1277
rect 259 -1286 263 -1236
rect 518 -1276 522 -1267
rect 591 -1276 595 -1219
rect 652 -1256 656 -1213
rect 828 -1228 832 -1219
rect 901 -1228 905 -1171
rect 962 -1208 966 -1165
rect 1310 -1189 1314 -1099
rect 1620 -1141 1624 -1099
rect 1721 -1165 1756 -1161
rect 1060 -1214 1082 -1210
rect 1411 -1213 1446 -1209
rect 828 -1232 905 -1228
rect 831 -1260 835 -1256
rect 750 -1264 835 -1260
rect 511 -1280 595 -1276
rect 158 -1290 263 -1286
rect 88 -1366 123 -1362
rect 259 -1399 263 -1290
rect 521 -1308 525 -1304
rect 472 -1312 525 -1308
rect 144 -1403 263 -1399
rect 271 -1363 296 -1359
rect 173 -1441 177 -1403
rect 271 -1409 275 -1363
rect 242 -1413 275 -1409
rect -91 -1445 177 -1441
rect -461 -1463 -250 -1459
rect 472 -1463 476 -1312
rect 521 -1416 525 -1312
rect 591 -1337 595 -1280
rect 606 -1337 610 -1328
rect 692 -1337 696 -1287
rect 591 -1341 696 -1337
rect 521 -1420 556 -1416
rect 692 -1444 696 -1341
rect 831 -1365 835 -1264
rect 901 -1289 905 -1232
rect 916 -1289 920 -1280
rect 1002 -1289 1006 -1239
rect 1277 -1276 1281 -1267
rect 1350 -1276 1354 -1219
rect 1411 -1256 1415 -1213
rect 1587 -1228 1591 -1219
rect 1660 -1228 1664 -1171
rect 1721 -1208 1725 -1165
rect 2046 -1189 2050 -1099
rect 2356 -1141 2360 -1099
rect 2457 -1165 2492 -1161
rect 1819 -1214 1837 -1210
rect 2147 -1213 2182 -1209
rect 1587 -1232 1664 -1228
rect 1590 -1260 1594 -1256
rect 1509 -1264 1594 -1260
rect 1277 -1280 1354 -1276
rect 901 -1293 1006 -1289
rect 831 -1369 866 -1365
rect 1002 -1402 1006 -1293
rect 1280 -1308 1284 -1304
rect 1241 -1312 1284 -1308
rect 887 -1406 1006 -1402
rect 1014 -1366 1039 -1362
rect 916 -1444 920 -1406
rect 1014 -1412 1018 -1366
rect 985 -1416 1018 -1412
rect 652 -1448 920 -1444
rect 1241 -1467 1245 -1312
rect 1280 -1416 1284 -1312
rect 1350 -1337 1354 -1280
rect 1365 -1337 1369 -1328
rect 1451 -1337 1455 -1287
rect 1350 -1341 1455 -1337
rect 1280 -1420 1315 -1416
rect 1451 -1443 1455 -1341
rect 1590 -1365 1594 -1264
rect 1660 -1289 1664 -1232
rect 1675 -1289 1679 -1280
rect 1761 -1289 1765 -1239
rect 2013 -1276 2017 -1267
rect 2086 -1276 2090 -1219
rect 2147 -1256 2151 -1213
rect 2323 -1228 2327 -1219
rect 2396 -1228 2400 -1171
rect 2457 -1208 2461 -1165
rect 2555 -1214 2571 -1210
rect 2323 -1232 2400 -1228
rect 2326 -1260 2330 -1256
rect 2245 -1264 2330 -1260
rect 2013 -1280 2090 -1276
rect 1660 -1293 1765 -1289
rect 1590 -1369 1625 -1365
rect 1761 -1402 1765 -1293
rect 2016 -1308 2020 -1304
rect 1965 -1312 2020 -1308
rect 1646 -1406 1765 -1402
rect 1773 -1366 1798 -1362
rect 1675 -1443 1679 -1406
rect 1773 -1412 1777 -1366
rect 1744 -1416 1777 -1412
rect 1406 -1447 1679 -1443
rect -469 -1480 -250 -1476
rect 1965 -1478 1969 -1312
rect 2016 -1416 2020 -1312
rect 2086 -1337 2090 -1280
rect 2101 -1337 2105 -1328
rect 2187 -1337 2191 -1287
rect 2086 -1341 2191 -1337
rect 2016 -1420 2051 -1416
rect 2187 -1443 2191 -1341
rect 2326 -1365 2330 -1264
rect 2396 -1289 2400 -1232
rect 2411 -1289 2415 -1280
rect 2497 -1289 2501 -1239
rect 2396 -1293 2501 -1289
rect 2326 -1369 2361 -1365
rect 2497 -1402 2501 -1293
rect 2382 -1406 2501 -1402
rect 2509 -1366 2534 -1362
rect 2411 -1443 2415 -1406
rect 2509 -1412 2513 -1366
rect 2480 -1416 2513 -1412
rect 2142 -1446 2415 -1443
rect -477 -1492 -250 -1488
rect -505 -1526 -482 -1522
rect -879 -1580 -591 -1576
rect -486 -1614 -482 -1526
rect -505 -1618 -482 -1614
rect -910 -1643 -600 -1639
rect -739 -1700 -593 -1696
rect -486 -1734 -482 -1618
rect -504 -1738 -482 -1734
rect -759 -1792 -593 -1788
rect -486 -1826 -482 -1738
rect -477 -1792 -473 -1692
rect -507 -1830 -482 -1826
rect -779 -1884 -593 -1880
rect -486 -1918 -482 -1830
rect -466 -1884 -462 -1667
rect -507 -1922 -482 -1918
rect -799 -1976 -593 -1972
rect -486 -2010 -482 -1922
rect -455 -1985 -451 -1642
rect -507 -2014 -482 -2010
rect -819 -2067 -591 -2063
rect -486 -2101 -482 -2014
rect -250 -2038 -234 -1642
rect -218 -2021 -202 -1667
rect -186 -2004 -170 -1692
rect -250 -2046 -213 -2038
rect -502 -2105 -482 -2101
rect -839 -2159 -591 -2155
rect -486 -2193 -482 -2105
rect -151 -2158 -135 -1709
rect -55 -1709 -51 -1653
rect -26 -1704 1184 -1696
rect -26 -1708 -17 -1704
rect -26 -1709 -22 -1708
rect -55 -1713 -22 -1709
rect 463 -1708 472 -1704
rect -26 -1755 -22 -1713
rect 463 -1755 467 -1708
rect 847 -1708 856 -1704
rect 847 -1755 851 -1708
rect 1180 -1733 1184 -1704
rect 1180 -1737 1266 -1733
rect 75 -1779 110 -1775
rect 564 -1779 599 -1775
rect 948 -1779 1017 -1775
rect 1262 -1779 1266 -1737
rect -59 -1842 -55 -1833
rect 14 -1842 18 -1785
rect 75 -1817 79 -1779
rect 75 -1822 102 -1817
rect -96 -1846 18 -1842
rect -505 -2197 -482 -2193
rect -859 -2251 -591 -2247
rect -486 -2285 -482 -2197
rect -505 -2289 -482 -2285
rect -119 -2284 -103 -1904
rect -96 -2219 -92 -1846
rect 14 -1903 18 -1846
rect 98 -1885 102 -1822
rect 430 -1842 434 -1833
rect 503 -1842 507 -1785
rect 564 -1822 568 -1779
rect 430 -1846 507 -1842
rect 814 -1842 818 -1833
rect 887 -1842 891 -1785
rect 948 -1822 952 -1779
rect 1363 -1803 1398 -1799
rect 814 -1846 891 -1842
rect 115 -1879 119 -1853
rect 115 -1883 123 -1879
rect 29 -1903 33 -1894
rect 115 -1903 119 -1883
rect 503 -1903 507 -1846
rect 604 -1879 608 -1853
rect 604 -1883 612 -1879
rect 518 -1903 522 -1894
rect 604 -1903 608 -1883
rect 887 -1903 891 -1846
rect 1022 -1879 1026 -1853
rect 1229 -1866 1233 -1857
rect 1302 -1866 1306 -1809
rect 1363 -1846 1367 -1803
rect 1229 -1870 1306 -1866
rect 1022 -1883 1030 -1879
rect 902 -1903 906 -1894
rect 1022 -1903 1026 -1883
rect 1302 -1903 1306 -1870
rect 1403 -1897 1407 -1877
rect 1464 -1897 1468 -1885
rect 14 -1907 1306 -1903
rect 98 -2130 106 -1918
rect 1302 -1927 1306 -1907
rect 1388 -1901 1468 -1897
rect 1317 -1927 1321 -1918
rect 1388 -1927 1393 -1901
rect 1302 -1931 1393 -1927
rect 199 -2075 205 -2005
rect 43 -2138 106 -2130
rect 43 -2151 47 -2138
rect 4 -2156 42 -2152
rect -96 -2223 -53 -2219
rect -1 -2230 5 -2156
rect -7 -2234 5 -2230
rect 13 -2199 44 -2195
rect -119 -2288 -43 -2284
rect 13 -2284 17 -2199
rect 54 -2236 58 -2228
rect 120 -2236 124 -2228
rect 191 -2236 195 -2204
rect -8 -2288 17 -2284
rect 28 -2240 195 -2236
rect -879 -2343 -591 -2339
rect -486 -2377 -482 -2289
rect -61 -2325 -57 -2288
rect 28 -2316 32 -2240
rect 191 -2314 195 -2240
rect 209 -2262 225 -1932
rect 243 -2123 247 -2076
rect 612 -2075 618 -2033
rect 234 -2128 242 -2124
rect 307 -2119 363 -2115
rect 234 -2215 238 -2128
rect 209 -2266 248 -2262
rect 242 -2302 246 -2266
rect 307 -2269 311 -2119
rect 477 -2162 481 -2089
rect 455 -2181 602 -2177
rect 317 -2212 321 -2198
rect 594 -2231 602 -2181
rect 594 -2236 608 -2231
rect 275 -2273 311 -2269
rect 322 -2256 381 -2252
rect 322 -2302 326 -2256
rect 503 -2272 532 -2268
rect 242 -2306 326 -2302
rect 28 -2320 50 -2316
rect 191 -2318 347 -2314
rect -61 -2329 36 -2325
rect 46 -2352 50 -2320
rect 155 -2324 183 -2320
rect 55 -2352 59 -2344
rect 121 -2352 125 -2344
rect -1 -2356 125 -2352
rect -505 -2381 -482 -2377
rect -932 -2570 -600 -2566
rect -739 -2627 -593 -2623
rect -486 -2661 -482 -2381
rect 0 -2556 4 -2356
rect 175 -2371 183 -2324
rect 175 -2376 250 -2371
rect 204 -2441 215 -2389
rect 242 -2513 250 -2376
rect 528 -2400 532 -2272
rect 624 -2290 640 -1960
rect 659 -2123 663 -2076
rect 650 -2128 658 -2124
rect 723 -2119 779 -2115
rect 650 -2243 654 -2128
rect 723 -2284 727 -2119
rect 733 -2240 737 -2198
rect 843 -2220 847 -2071
rect 1056 -2075 1062 -2058
rect 867 -2208 1052 -2203
rect 1068 -2259 1072 -1988
rect 1103 -2123 1107 -2076
rect 1094 -2128 1102 -2124
rect 1173 -2119 1229 -2115
rect 1094 -2215 1098 -2128
rect 1068 -2263 1107 -2259
rect 1173 -2257 1177 -2119
rect 1183 -2212 1187 -2198
rect 1292 -2199 1296 -2076
rect 1134 -2261 1177 -2257
rect 1188 -2256 1247 -2252
rect 684 -2288 727 -2284
rect 738 -2284 797 -2280
rect 624 -2294 657 -2290
rect 640 -2330 644 -2294
rect 738 -2330 742 -2284
rect 903 -2300 932 -2296
rect 640 -2334 742 -2330
rect 258 -2408 532 -2400
rect 258 -2504 266 -2408
rect 924 -2416 932 -2300
rect 1068 -2302 1072 -2263
rect 1188 -2302 1192 -2256
rect 1353 -2272 1382 -2268
rect 1068 -2306 1192 -2302
rect 1032 -2335 1058 -2331
rect 272 -2424 932 -2416
rect 272 -2495 280 -2424
rect 1374 -2432 1382 -2272
rect 1388 -2336 1393 -1931
rect 284 -2440 1382 -2432
rect 284 -2490 292 -2440
rect 272 -2499 292 -2495
rect 258 -2508 292 -2504
rect 242 -2517 292 -2513
rect -504 -2665 -482 -2661
rect -759 -2719 -593 -2715
rect -486 -2753 -482 -2665
rect -507 -2757 -482 -2753
rect -779 -2811 -593 -2807
rect -486 -2845 -482 -2757
rect -507 -2849 -482 -2845
rect -799 -2903 -593 -2899
rect -486 -2937 -482 -2849
rect -507 -2941 -482 -2937
rect -819 -2994 -591 -2990
rect -486 -3028 -482 -2941
rect -125 -2798 -91 -2794
rect -125 -2999 -121 -2798
rect -6 -2824 18 -2820
rect -472 -3003 -121 -2999
rect -115 -2891 -91 -2887
rect -502 -3032 -482 -3028
rect -839 -3086 -591 -3082
rect -486 -3120 -482 -3032
rect -115 -3091 -111 -2891
rect 14 -2913 18 -2824
rect -6 -2917 18 -2913
rect -472 -3095 -111 -3091
rect -105 -2983 -91 -2979
rect -505 -3124 -482 -3120
rect -859 -3178 -591 -3174
rect -486 -3212 -482 -3124
rect -105 -3186 -101 -2983
rect 14 -3005 18 -2917
rect -6 -3009 18 -3005
rect -472 -3190 -101 -3186
rect -505 -3216 -482 -3212
rect -879 -3270 -591 -3266
rect -486 -3304 -482 -3216
rect -95 -3275 -91 -3072
rect 14 -3098 18 -3009
rect -6 -3102 18 -3098
rect -472 -3279 -91 -3275
rect 14 -3304 18 -3102
rect -505 -3308 18 -3304
<< m3contact >>
rect -537 -73 -532 -68
<< m123contact >>
rect -896 163 -891 168
rect -722 163 -717 168
rect -643 163 -638 168
rect -654 154 -649 159
rect -879 54 -874 59
rect -538 106 -533 111
rect -731 82 -726 87
rect -643 82 -638 87
rect -722 54 -717 59
rect -664 54 -659 59
rect -731 -27 -726 -22
rect -643 -27 -638 -22
rect -593 -101 -588 -96
rect -593 -192 -588 -187
rect -593 -284 -588 -279
rect -593 -376 -588 -371
rect -591 -468 -586 -463
rect -591 -559 -586 -554
rect -591 -651 -586 -646
rect -400 -213 -395 -208
rect -426 -232 -421 -227
rect -440 -249 -435 -244
rect -453 -439 -448 -434
rect 2 -120 7 -115
rect 746 -120 751 -115
rect 1515 -120 1520 -115
rect 2249 -120 2254 -115
rect -243 -213 -238 -208
rect -243 -232 -238 -227
rect -243 -249 -238 -244
rect 3 -394 8 -389
rect -277 -439 -272 -434
rect 746 -397 751 -392
rect 1530 -397 1535 -392
rect 2266 -397 2271 -392
rect -591 -743 -586 -738
rect -630 -888 -625 -883
rect -593 -894 -588 -889
rect -593 -985 -588 -980
rect -593 -1077 -588 -1072
rect -593 -1169 -588 -1164
rect -591 -1261 -586 -1256
rect -591 -1352 -586 -1347
rect -591 -1444 -586 -1439
rect -400 -1006 -395 -1001
rect -426 -1025 -421 -1020
rect -440 -1042 -435 -1037
rect -453 -1232 -448 -1227
rect 31 -913 36 -908
rect 775 -913 780 -908
rect 1544 -913 1549 -908
rect 2278 -913 2283 -908
rect -214 -1006 -209 -1001
rect -214 -1025 -209 -1020
rect -214 -1042 -209 -1037
rect 32 -1187 37 -1182
rect -248 -1232 -243 -1227
rect 775 -1190 780 -1185
rect 1559 -1190 1564 -1185
rect 2295 -1190 2300 -1185
rect -591 -1536 -586 -1531
rect -593 -1657 -588 -1652
rect -593 -1748 -588 -1743
rect -593 -1840 -588 -1835
rect -593 -1932 -588 -1927
rect -591 -2024 -586 -2019
rect -591 -2115 -586 -2110
rect -591 -2207 -586 -2202
rect 287 -1832 295 -1827
rect 703 -1832 708 -1827
rect 1153 -1832 1161 -1827
rect 1493 -1853 1498 -1848
rect -591 -2299 -586 -2294
rect 387 -2131 392 -2126
rect 405 -2268 410 -2263
rect -593 -2584 -588 -2579
rect 519 -2336 524 -2331
rect 803 -2131 808 -2126
rect 1253 -2131 1258 -2126
rect 821 -2296 826 -2291
rect 937 -2297 942 -2292
rect 545 -2348 550 -2343
rect 663 -2345 668 -2340
rect 537 -2374 542 -2369
rect 1271 -2268 1276 -2263
rect 954 -2309 959 -2304
rect 943 -2328 948 -2323
rect 1048 -2345 1053 -2340
rect 1430 -2289 1435 -2284
rect 1430 -2305 1435 -2300
rect 1430 -2314 1435 -2309
rect 1430 -2323 1435 -2318
rect -593 -2675 -588 -2670
rect -593 -2767 -588 -2762
rect -593 -2859 -588 -2854
rect -591 -2951 -586 -2946
rect -591 -3042 -586 -3037
rect -591 -3134 -586 -3129
rect -591 -3226 -586 -3221
<< metal3 >>
rect -912 163 -896 167
rect -717 163 -643 167
rect -912 66 -908 163
rect -653 86 -649 154
rect -726 82 -643 86
rect -912 58 -907 66
rect -912 54 -879 58
rect -717 54 -664 58
rect -912 -97 -907 54
rect -653 -23 -649 82
rect -726 -27 -643 -23
rect -537 -68 -533 106
rect -912 -101 -593 -97
rect -616 -188 -612 -101
rect -616 -192 -593 -188
rect -616 -280 -612 -192
rect -395 -213 -243 -209
rect -421 -232 -243 -228
rect -435 -249 -243 -245
rect -616 -284 -593 -280
rect -616 -372 -612 -284
rect -616 -376 -593 -372
rect -616 -464 -612 -376
rect 3 -389 7 -120
rect 746 -392 750 -120
rect 1516 -393 1520 -120
rect 1516 -397 1530 -393
rect 2250 -393 2254 -120
rect 2250 -397 2266 -393
rect -448 -439 -277 -435
rect -616 -468 -591 -464
rect -616 -555 -612 -468
rect -616 -559 -591 -555
rect -616 -647 -612 -559
rect -616 -651 -591 -647
rect -616 -739 -612 -651
rect -616 -743 -591 -739
rect -616 -890 -612 -743
rect -616 -894 -593 -890
rect -616 -981 -612 -894
rect -616 -985 -593 -981
rect -616 -1073 -612 -985
rect -395 -1006 -214 -1002
rect -421 -1025 -214 -1021
rect -435 -1042 -214 -1038
rect -616 -1077 -593 -1073
rect -616 -1165 -612 -1077
rect -616 -1169 -593 -1165
rect -616 -1257 -612 -1169
rect 32 -1182 36 -913
rect 775 -1185 779 -913
rect 1545 -1186 1549 -913
rect 1545 -1190 1559 -1186
rect 2279 -1186 2283 -913
rect 2279 -1190 2295 -1186
rect -448 -1232 -248 -1228
rect -616 -1261 -591 -1257
rect -616 -1348 -612 -1261
rect -616 -1352 -591 -1348
rect -616 -1440 -612 -1352
rect -616 -1444 -591 -1440
rect -616 -1532 -612 -1444
rect -616 -1536 -591 -1532
rect -616 -1653 -612 -1536
rect -616 -1657 -593 -1653
rect -616 -1744 -612 -1657
rect -616 -1748 -593 -1744
rect -616 -1836 -612 -1748
rect -616 -1840 -593 -1836
rect -616 -1928 -612 -1840
rect -616 -1932 -593 -1928
rect -616 -2020 -612 -1932
rect -616 -2024 -591 -2020
rect -616 -2111 -612 -2024
rect -616 -2115 -591 -2111
rect -616 -2203 -612 -2115
rect 287 -2127 295 -1832
rect 703 -1895 707 -1832
rect 612 -1899 707 -1895
rect 612 -1946 616 -1899
rect 519 -1950 616 -1946
rect 287 -2131 387 -2127
rect -616 -2207 -591 -2203
rect -616 -2295 -612 -2207
rect 287 -2264 295 -2131
rect 287 -2268 405 -2264
rect -616 -2299 -591 -2295
rect -616 -2580 -612 -2299
rect 287 -2344 295 -2268
rect 519 -2331 523 -1950
rect 1153 -1968 1161 -1832
rect 1493 -1927 1497 -1853
rect 937 -1976 1161 -1968
rect 1401 -1931 1497 -1927
rect 703 -2131 803 -2127
rect 703 -2292 711 -2131
rect 703 -2296 821 -2292
rect 937 -2292 941 -1976
rect 1153 -2131 1253 -2127
rect 1153 -2264 1161 -2131
rect 1153 -2268 1271 -2264
rect 703 -2340 711 -2296
rect 287 -2348 545 -2344
rect 668 -2345 711 -2340
rect 287 -2384 295 -2348
rect 703 -2356 711 -2345
rect 935 -2309 954 -2305
rect 935 -2356 939 -2309
rect 703 -2364 939 -2356
rect 943 -2360 948 -2328
rect 1153 -2341 1161 -2268
rect 1401 -2285 1405 -1931
rect 1401 -2289 1430 -2285
rect 1053 -2345 1161 -2341
rect 1402 -2305 1430 -2301
rect 1402 -2360 1406 -2305
rect 943 -2368 1406 -2360
rect 1414 -2314 1430 -2310
rect 1414 -2372 1418 -2314
rect 542 -2374 1418 -2372
rect 538 -2380 1418 -2374
rect 1426 -2384 1430 -2319
rect 287 -2392 1430 -2384
rect -616 -2584 -593 -2580
rect -616 -2671 -612 -2584
rect -616 -2675 -593 -2671
rect -616 -2763 -612 -2675
rect -616 -2767 -593 -2763
rect -616 -2855 -612 -2767
rect -616 -2859 -593 -2855
rect -616 -2947 -612 -2859
rect -616 -2951 -591 -2947
rect -616 -3038 -612 -2951
rect -616 -3042 -591 -3038
rect -616 -3130 -612 -3042
rect -616 -3134 -591 -3130
rect -616 -3222 -612 -3134
rect -616 -3226 -591 -3222
<< labels >>
rlabel metal1 -719 3 -717 4 1 D2
rlabel metal1 -718 113 -716 114 1 D0
rlabel metal1 -888 120 -884 123 1 S0
rlabel metal1 -880 165 -878 166 4 VDD
rlabel metal1 -880 83 -878 84 2 GND
rlabel metal1 -862 117 -858 118 1 S0comp
rlabel metal1 -814 108 -810 109 1 S0comp
rlabel metal2 -824 120 -821 122 1 S1comp
rlabel metal1 -885 11 -881 13 1 S1
rlabel metal1 -858 8 -855 9 1 S1comp
rlabel metal1 -814 -1 -810 0 1 S0comp
rlabel metal1 -812 12 -808 14 1 S1
rlabel metal1 -645 0 -641 1 1 S0
rlabel metal2 -647 12 -644 13 1 S1
rlabel metal1 -552 3 -549 4 7 D3
rlabel metal1 -641 109 -637 110 1 S0
rlabel metal2 -647 121 -644 122 1 S1comp
rlabel metal1 -547 112 -544 113 7 D1
rlabel metal2 -230 -132 -226 -131 1 GND
rlabel metal1 595 -114 598 -113 1 B1new
rlabel metal1 1474 -114 1477 -113 1 B2new
rlabel metal1 3 -114 6 -113 1 B0new
rlabel metal1 2240 -114 2243 -113 1 B3new
rlabel metal1 -496 -152 -493 -151 1 A3_add
rlabel metal1 -497 -244 -494 -243 1 A2_add
rlabel metal1 -498 -336 -495 -335 1 A1_add
rlabel metal1 -496 -438 -493 -437 1 A0_add
rlabel metal1 -496 -519 -493 -518 1 B3_add
rlabel metal1 -498 -611 -495 -610 1 B2_add
rlabel metal1 -500 -706 -497 -705 1 B1_add
rlabel metal1 -499 -795 -496 -794 1 B0_add
rlabel metal1 -747 -114 -745 -112 1 A3
rlabel metal1 -767 -114 -765 -112 1 A2
rlabel metal1 -787 -114 -785 -112 1 A1
rlabel metal1 -807 -114 -805 -112 1 A0
rlabel metal1 -827 -114 -825 -112 1 B3
rlabel metal1 -847 -114 -845 -112 1 B2
rlabel metal1 -867 -114 -865 -112 1 B1
rlabel metal1 -887 -114 -885 -112 1 B0
rlabel metal3 -615 -101 -612 -99 5 VDD
rlabel metal1 -668 -85 -664 -82 1 D0
rlabel metal2 -398 12 -396 13 1 k
rlabel metal2 301 -417 304 -416 1 sum0
rlabel metal2 1043 -421 1047 -419 1 sum1
rlabel metal2 1804 -420 1807 -419 1 sum2
rlabel metal2 2538 -420 2542 -418 1 sum3
rlabel metal1 2596 -567 2598 -566 1 final_carry
rlabel metal2 -201 -925 -197 -924 1 GND
rlabel metal1 -352 -807 -347 -805 1 D1
rlabel metal1 32 -907 35 -905 1 B0new_sub
rlabel metal1 624 -907 628 -906 1 B1new_sub
rlabel metal1 1503 -907 1507 -906 1 B2new_sub
rlabel metal1 2269 -907 2273 -906 1 B3new_sub
rlabel metal2 330 -1210 333 -1209 1 diff0
rlabel metal2 1074 -1213 1076 -1212 1 diff1
rlabel metal2 1833 -1213 1836 -1212 1 diff2
rlabel metal2 2567 -1213 2569 -1212 1 diff3
rlabel metal1 2625 -1360 2627 -1359 1 final_borrow
rlabel metal1 -499 -1588 -496 -1587 1 B0_sub
rlabel metal1 -500 -1499 -497 -1498 1 B1_sub
rlabel metal1 -499 -1404 -495 -1403 1 B2_sub
rlabel metal1 -496 -1312 -492 -1311 1 B3_sub
rlabel metal1 -496 -1231 -494 -1230 1 A0_sub
rlabel metal1 -500 -1129 -497 -1128 1 A1_sub
rlabel metal1 -499 -1037 -496 -1036 1 A2_sub
rlabel metal1 -497 -945 -492 -944 1 A3_sub
rlabel metal1 -496 -1708 -493 -1707 1 A3_comp
rlabel metal1 -497 -1800 -494 -1799 1 A2_comp
rlabel metal1 -498 -1892 -495 -1891 1 A1_comp
rlabel metal1 -496 -1994 -493 -1993 1 A0_comp
rlabel metal1 -496 -2075 -493 -2074 1 B3_comp
rlabel metal1 -498 -2167 -495 -2166 1 B2_comp
rlabel metal1 -498 -2262 -495 -2261 1 B1_comp
rlabel metal1 -499 -2351 -496 -2350 1 B0_comp
rlabel metal2 712 -2287 715 -2286 1 B1comp
rlabel metal1 453 -2507 455 -2506 1 lesser
rlabel metal1 300 -2516 302 -2515 1 L3
rlabel metal1 300 -2507 302 -2506 1 L2
rlabel metal1 300 -2498 302 -2497 1 L1
rlabel metal1 300 -2489 302 -2488 1 L0
rlabel metal1 182 -2492 184 -2491 1 greater
rlabel metal1 33 -2489 35 -2488 1 G0
rlabel metal1 33 -2497 35 -2496 1 G1
rlabel metal1 33 -2505 35 -2504 1 G2
rlabel metal1 33 -2513 35 -2512 1 G3
rlabel metal3 290 -2360 293 -2358 1 E3
rlabel metal1 257 -1831 259 -1830 1 E3
rlabel metal2 178 -2360 180 -2359 1 L3
rlabel metal1 460 -2134 463 -2133 1 G2
rlabel metal1 478 -2271 481 -2270 1 L2
rlabel metal1 690 -2175 695 -2173 1 A1comp
rlabel metal1 876 -2134 879 -2133 1 G1
rlabel metal1 699 -1831 701 -1830 1 E2
rlabel metal1 894 -2299 897 -2298 1 L1
rlabel metal1 161 -2360 163 -2359 1 G3
rlabel metal2 1162 -2261 1166 -2259 1 B0comp
rlabel metal1 1488 -1851 1491 -1850 1 E0
rlabel metal3 1427 -2326 1430 -2325 1 E3
rlabel metal3 1424 -2304 1427 -2303 1 E1
rlabel metal3 1424 -2288 1427 -2287 1 E0
rlabel metal1 1579 -2313 1581 -2311 7 equal
rlabel metal1 1117 -1831 1119 -1830 1 E1
rlabel metal2 1377 -2359 1380 -2357 1 L0
rlabel metal1 1360 -2359 1363 -2357 1 G0
rlabel metal1 1326 -2134 1329 -2133 1 G0
rlabel metal1 1344 -2271 1347 -2270 1 L0
rlabel metal3 1424 -2313 1427 -2312 1 E2
rlabel metal1 910 -2355 913 -2354 1 G1
rlabel metal2 927 -2354 930 -2353 1 L1
rlabel metal3 699 -2343 702 -2342 1 E3.E2
rlabel metal3 1065 -2344 1068 -2343 1 E3.E2.E1
rlabel metal1 275 -2175 278 -2174 1 A2comp
rlabel metal2 297 -2272 299 -2271 1 B2comp
rlabel metal1 -16 -2194 -13 -2193 1 A3comp
rlabel metal1 -496 -2635 -493 -2634 1 A3_and
rlabel metal1 -497 -2727 -492 -2726 1 A2_and
rlabel metal1 -498 -2819 -495 -2818 1 A1_and
rlabel metal1 -496 -3002 -493 -3001 1 B3_and
rlabel metal1 -498 -3094 -495 -3093 1 B2_and
rlabel metal1 -498 -3189 -495 -3188 1 B1_and
rlabel metal1 -499 -3278 -496 -3277 1 B0_and
rlabel metal1 -496 -2911 -493 -2910 1 A0_and
rlabel metal1 2 -2794 4 -2793 1 Ans3
rlabel metal1 2 -2887 4 -2886 1 Ans2
rlabel metal1 2 -2979 4 -2978 1 Ans1
rlabel metal1 2 -3072 4 -3071 1 Ans0
<< end >>
