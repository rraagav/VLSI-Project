magic
tech scmos
timestamp 1700487792
<< nwell >>
rect -2 0 58 24
<< ntransistor >>
rect 10 -37 14 -29
rect 31 -37 35 -29
<< ptransistor >>
rect 10 8 14 16
rect 31 8 35 16
<< ndiffusion >>
rect 4 -31 10 -29
rect 4 -35 5 -31
rect 9 -35 10 -31
rect 4 -37 10 -35
rect 14 -37 31 -29
rect 35 -31 52 -29
rect 35 -35 38 -31
rect 42 -35 52 -31
rect 35 -37 52 -35
<< pdiffusion >>
rect 4 14 10 16
rect 4 10 5 14
rect 9 10 10 14
rect 4 8 10 10
rect 14 14 31 16
rect 14 10 15 14
rect 19 10 31 14
rect 14 8 31 10
rect 35 14 52 16
rect 35 10 38 14
rect 42 10 52 14
rect 35 8 52 10
<< ndcontact >>
rect 5 -35 9 -31
rect 38 -35 42 -31
<< pdcontact >>
rect 5 10 9 14
rect 15 10 19 14
rect 38 10 42 14
<< polysilicon >>
rect 10 16 14 19
rect 31 16 35 19
rect 10 -29 14 8
rect 31 -29 35 8
rect 10 -40 14 -37
rect 31 -45 35 -37
<< polycontact >>
rect 6 -11 10 -7
rect 27 -23 31 -19
<< metal1 >>
rect -2 32 46 36
rect 5 14 9 32
rect 38 14 42 32
rect 2 -11 6 -7
rect 15 -11 19 10
rect 15 -15 58 -11
rect 2 -23 27 -19
rect 38 -31 42 -15
rect 5 -45 9 -35
rect -2 -49 16 -45
<< labels >>
rlabel metal1 2 34 4 35 4 VDD
rlabel metal1 2 -48 4 -47 2 GND
rlabel metal1 51 -14 54 -13 1 Vout
rlabel metal1 3 -10 5 -9 1 VA
rlabel metal1 3 -22 5 -21 1 VB
<< end >>
