* SPICE3 file created from xnor.ext - technology: scmos
.include TSMC_180nm.txt

.param SUPPLY = 1.8
.param LAMBDA = 0.18u
.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}
.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd VDD gnd 'Supply'

Vin_A VA gnd DC(0)
Vin_B VB gnd DC(0)

.option scale=0.09u

M1000 a_266_9# VB a_266_n36# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=136 ps=50
M1001 a_440_n11# a_339_57# VDD w_424_n19# CMOSP w=8 l=4
+  ad=136 pd=50 as=784 ps=340
M1002 VDD a_266_9# a_339_57# w_323_49# CMOSP w=8 l=4
+  ad=0 pd=0 as=136 ps=50
M1003 a_339_57# a_266_9# a_339_12# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=136 ps=50
M1004 VDD a_354_n52# a_440_n11# w_424_n19# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1005 Vout a_440_n11# VDD w_492_n19# CMOSP w=8 l=4
+  ad=48 pd=28 as=0 ps=0
M1006 a_354_n97# a_266_9# GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=240 ps=140
M1007 a_266_9# VA VDD w_250_1# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1008 a_354_n52# VB a_354_n97# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1009 a_339_57# VA VDD w_323_49# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1010 a_339_12# VA GND Gnd CMOSN w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1011 a_440_n56# a_339_57# GND Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1012 VDD VB a_266_9# w_250_1# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1013 a_354_n52# a_266_9# VDD w_338_n60# CMOSP w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1014 a_440_n11# a_354_n52# a_440_n56# Gnd CMOSN w=8 l=4
+  ad=136 pd=50 as=0 ps=0
M1015 a_266_n36# VA GND Gnd CMOSN w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1016 VDD VB a_354_n52# w_338_n60# CMOSP w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1017 Vout a_440_n11# GND Gnd CMOSN w=8 l=4
+  ad=48 pd=28 as=0 ps=0
C0 a_266_9# GND 0.26fF
C1 w_338_n60# a_354_n52# 0.03fF
C2 w_492_n19# a_440_n11# 0.11fF
C3 a_266_9# VDD 0.03fF
C4 VA a_339_57# 0.03fF
C5 w_338_n60# VB 0.11fF
C6 w_492_n19# VDD 0.03fF
C7 w_338_n60# a_266_9# 0.11fF
C8 w_424_n19# a_339_57# 0.11fF
C9 w_250_1# VB 0.11fF
C10 w_250_1# a_266_9# 0.03fF
C11 w_323_49# VDD 0.05fF
C12 a_440_n11# Vout 0.03fF
C13 GND Vout 0.03fF
C14 a_339_57# a_440_n11# 0.03fF
C15 VDD Vout 0.03fF
C16 VB a_354_n52# 0.10fF
C17 a_266_9# a_354_n52# 0.03fF
C18 VDD a_339_57# 0.11fF
C19 w_424_n19# a_440_n11# 0.03fF
C20 a_266_9# VB 0.10fF
C21 VA VDD 0.09fF
C22 w_424_n19# VDD 0.05fF
C23 w_250_1# VA 0.11fF
C24 w_323_49# a_266_9# 0.11fF
C25 VDD a_440_n11# 0.03fF
C26 w_492_n19# Vout 0.03fF
C27 a_266_9# a_339_57# 0.10fF
C28 w_424_n19# a_354_n52# 0.11fF
C29 VA a_266_9# 0.03fF
C30 w_338_n60# VDD 0.05fF
C31 w_250_1# VDD 0.05fF
C32 w_323_49# a_339_57# 0.03fF
C33 w_323_49# VA 0.11fF
C34 a_354_n52# a_440_n11# 0.10fF
C35 GND a_354_n52# 0.09fF
C36 VDD a_354_n52# 0.03fF
C37 VB GND 0.17fF
C38 Vout Gnd 0.10fF
C39 a_440_n11# Gnd 0.51fF
C40 a_354_n52# Gnd 0.76fF
C41 GND Gnd 4.98fF
C42 VB Gnd 1.33fF
C43 a_339_57# Gnd 0.88fF
C44 VDD Gnd 0.04fF
C45 a_266_9# Gnd 1.29fF
C46 VA Gnd 1.31fF
C47 w_338_n60# Gnd 1.45fF
C48 w_492_n19# Gnd 0.67fF
C49 w_424_n19# Gnd 1.45fF
C50 w_250_1# Gnd 0.31fF
C51 w_323_49# Gnd 1.45fF

.tran 1n 800n
.control
run
plot v(VA) v(VB)+2 v(Vout)+4
.end
.endc