magic
tech scmos
timestamp 1699268865
<< nwell >>
rect -2 0 26 24
<< ntransistor >>
rect 10 -31 14 -23
<< ptransistor >>
rect 10 8 14 16
<< ndiffusion >>
rect 4 -25 10 -23
rect 4 -29 5 -25
rect 9 -29 10 -25
rect 4 -31 10 -29
rect 14 -25 20 -23
rect 14 -29 15 -25
rect 19 -29 20 -25
rect 14 -31 20 -29
<< pdiffusion >>
rect 4 14 10 16
rect 4 10 5 14
rect 9 10 10 14
rect 4 8 10 10
rect 14 14 20 16
rect 14 10 15 14
rect 19 10 20 14
rect 14 8 20 10
<< ndcontact >>
rect 5 -29 9 -25
rect 15 -29 19 -25
<< pdcontact >>
rect 5 10 9 14
rect 15 10 19 14
<< polysilicon >>
rect 10 16 14 19
rect 10 -23 14 8
rect 10 -34 14 -31
<< polycontact >>
rect 6 -11 10 -7
<< metal1 >>
rect -2 32 26 36
rect 5 14 9 32
rect 2 -11 6 -7
rect 15 -11 19 10
rect 15 -15 27 -11
rect 15 -25 19 -15
rect 5 -39 9 -29
rect -2 -43 26 -39
<< labels >>
rlabel metal1 3 -10 5 -9 1 Vin
rlabel metal1 19 -14 21 -13 1 Vout
rlabel metal1 2 34 4 35 4 VDD
rlabel metal1 2 -42 4 -41 2 GND
<< end >>
